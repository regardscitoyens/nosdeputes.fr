Parlementaire:
  depute_1001:
    fonctions:
      - délégation chargée de la communication audiovisuelle et de la presse / président / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1001
    adresses:
      - Hôtel de Ville BP 19 59831 Lambersart cedex Téléphone : 03 20 08 44 44 Télécopie : 03 20 08 44 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 53 Télécopie : 01 40 63 79 37 
    circonscription: Nord (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Daubresse
    place_hemicycle: 346
    autresmandats:
      - Maire de Lambersart, Nord (28129 habitants)
    mails:
      - mpdaubresse@ville-lambersart.fr
      - mpdaubresse@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1001.asp
    profession: Ancien directeur d'une société de recrutement
    site_web: http://www.mpdaubresse.com
    debut_mandat: 20/06/2007
    nom: Marc-Philippe Daubresse
    type: depute
  depute_1012:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 1012
    extras:
      - haut conseil du secteur public / membre titulaire
      - conseil d'orientation de la simplification administrative / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 4 Rue du Docteur Mehier BP 49 01152 Lagnieu Cedex Téléphone : 04 74 35 13 58  Télécopie : 04 74 35 74 93 
    circonscription: Ain (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Verpillière
    place_hemicycle: 40
    autresmandats:
      - Membre du conseil général (Ain)
    mails:
      - cdelaverpilliere@assemblee-nationale.fr
      - charlesdelaverpilliere@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1012.asp
    profession: Conseiller d'Etat
    site_web: http://www.charlesdelaverpilliere.com
    debut_mandat: 20/06/2007
    nom: Charles de La Verpillière
    type: depute
  depute_1020:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 1020
    extras:
      - comité consultatif national d'Éthique pour les sciences de la vie et de la santé / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (15ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bernard Debré
    place_hemicycle: 10
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Conseiller de Paris
    mails:
      - bdebre@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1020.asp
    profession: Chirurgien des hôpitaux, professeur des Universités
    site_web: http://www.bernarddebre.fr
    debut_mandat: 20/06/2007
    nom: Bernard Debré
    type: depute
  depute_1029:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1029
    adresses:
      - 4 Rue Chaulan 13400 Aubagne Téléphone : 04 42 82 20 10 Télécopie : 04 42 82 20 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Deflesselles
    place_hemicycle: 253
    autresmandats:
      - Membre du conseil régional (Provence-Alpes-Côte-d'Azur)
    mails:
      - bdeflesselles@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1029.asp
    profession: Ingénieur
    site_web: http://www.bernarddeflesselles.com
    debut_mandat: 20/06/2007
    nom: Bernard Deflesselles
    type: depute
  depute_1031:
    place_hemicycle: 52
    fonctions:
      - commission des affaires européennes / membre / 
      - commission chargée de l'application de l'article 26 de la constitution / secrétaire / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Maire de Courtieux, Oise (172 habitants)
      - Membre du conseil général (Oise)
      - Président de la communauté de communes du canton d'Attichy
    sexe: H
    id_an: 1031
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1031.asp
    mails:
      - ldegauchy@assemblee-nationale.fr
    adresses:
      - Rue d'Angoulême 60350 Courtieux Téléphone : 03 44 42 19 78 Télécopie : 03 44 42 90 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Horticulteur
    debut_mandat: 20/06/2007
    nom_de_famille: Degauchy
    nom: Lucien Degauchy
    type: depute
  depute_1032:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 1032
    adresses:
      - Permanence parlementaire 7 Bis Place de la Cité 24000 Périgueux Téléphone : 05 53 46 72 45 Télécopie : 05 53 09 08 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 73 35 Télécopie : 01 40 63 78 98 
    circonscription: Dordogne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Deguilhem
    place_hemicycle: 638
    autresmandats:
      - Membre du Conseil municipal de Saint-Aquilin, Dordogne (452 habitants)
      - Membre du conseil général (Dordogne)
    mails:
      - pascaldeguilhem@free.fr
      - pdeguilhem@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1032.asp
    profession: Professeur d'Education physique (Université Bordeaux IV)
    site_web: http://pascaldeguilhem.free.fr
    debut_mandat: 20/06/2007
    nom: Pascal Deguilhem
    type: depute
  depute_1048:
    place_hemicycle: 533
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Maire de Dunkerque, Nord (70776 habitants)
    sexe: H
    id_an: 1048
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1048.asp
    mails:
      - mdelebarre@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville BP 6537 59386 Dunkerque cedex 1 Téléphone : 03 28 26 26 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (13ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Préfet
    debut_mandat: 20/06/2007
    nom_de_famille: Delebarre
    nom: Michel Delebarre
    type: depute
  depute_1058:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 1058
    extras:
      - conseil national de la sécurité routière / membre titulaire
    adresses:
      - Hôtel de Ville BP 141 94321 Thiais cedex Téléphone : 01 48 92 42 01 Télécopie : 01 48 53 47 20 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Dell'Agnola
    place_hemicycle: 357
    autresmandats:
      - Maire de Thiais, Val-de-Marne (28244 habitants)
    mails:
      - rdellagnola@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1058.asp
    profession: Attaché principal d'administration au ministère de la justice
    site_web: http://www.richard-dellagnola.com
    debut_mandat: 20/06/2007
    nom: Richard Dell'Agnola
    type: depute
  depute_1066:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 1066
    adresses:
      - Assemblée nationale 126 Rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville Avenue de la Côte d'Argent 33470 Le Teich Téléphone : 05 56 22 33 66 Télécopie : 05 56 22 83 24 
    circonscription: Gironde (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Deluga
    place_hemicycle: 404
    autresmandats:
      - Vice-président de la communauté d'agglomération du Bassin d'Arcachon sud
      - Maire du Teich, Gironde (4822 habitants)
    mails:
      - f.deluga@leteich.fr
      - fdeluga@assemblee-nationale.fr
      - contact@francoisdeluga.net
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1066.asp
    profession: Agent général d'assurances
    site_web: http://www.francoisdeluga.net
    debut_mandat: 01/12/2008
    nom: François Deluga
    type: depute
  depute_1079:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 1079
    extras:
      - conseil supérieur de l'énergie / membre titulaire
      - conseil de l'immobilier de l'etat / membre titulaire
    adresses:
      - Secrétariat parlementaire 19 Rue des Granges 61000 Alençon Téléphone : 02 33 32 09 53 Télécopie : 02 33 26 97 10 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Orne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Deniaud
    place_hemicycle: 100
    autresmandats:
      - Membre du conseil régional (Basse Normandie)
    mails:
      - ydeniaud@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1079.asp
    profession: Cadre commercial
    site_web: http://www.yves-deniaud.org
    debut_mandat: 20/06/2007
    nom: Yves Deniaud
    type: depute
  depute_1085:
    place_hemicycle: 21
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 1085
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1085.asp
    mails:
      - bernarddepierre@wanadoo.fr
      - bdepierre@assemblee-nationale.fr
    adresses:
      - Permanence 17 Rue Diderot 21000 Dijon Téléphone : 03 80 73 34 47 Télécopie : 03 80 72 28 56 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côte-d'Or (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.bernard-depierre.com
    profession: Consultant 
    debut_mandat: 20/06/2007
    nom_de_famille: Depierre
    nom: Bernard Depierre
    type: depute
  depute_1092:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des lois / membre / 
    sexe: H
    id_an: 1092
    extras:
      - conseil d'orientation de l'observatoire de l'emploi public / membre titulaire
      - conseil d'orientation de la simplification administrative / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 51 Rue Gustave Delory 59047 Lille cedex Téléphone : 03 59 73 66 90 
    circonscription: Nord (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Derosier
    place_hemicycle: 528
    autresmandats:
      - Président du conseil général (Nord)
    mails:
      - bderosier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1092.asp
    profession: Instituteur retraité
    debut_mandat: 20/06/2007
    nom: Bernard Derosier
    type: depute
  depute_1094:
    fonctions:
      - commission des affaires européennes / secrétaire / 
      - délégation chargée des activités internationales / membre / 
      - assemblée nationale / secrétaire / 27/06/2007
      - délégation chargée des représentants d'intérêts / membre / 
      - délégation spéciale chargée de la question des groupes d'intérêt / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1094
    adresses:
      - Hôtel de Ville 02700 Tergnier Téléphone : 03 23 57 11 27 Télécopie : 03 23 57 65 95 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 4 Avenue de Compiègne 02200 Soissons Téléphone : 03 23 59 05 41 Télécopie : 03 23 59 53 12 
    circonscription: Aisne (4ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Desallangre
    place_hemicycle: 581
    autresmandats:
      - Maire de Tergnier, Aisne (15069 habitants)
      - Président de la communauté de communes Chaugny Tergnier
    mails:
      - jdesallangre@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1094.asp
    profession: Journaliste
    site_web: http://www.jacques-desallangre.org/accueil.php
    debut_mandat: 20/06/2007
    nom: Jacques Desallangre
    type: depute
  depute_1116:
    fonctions:
      - commission des affaires étrangères / vice-président / 
    sexe: H
    id_an: 1116
    adresses:
      - Hôtel de Ville,  11 Boulevard Jean Pain BP 1066 38021 Grenoble cedex 1 Téléphone : 04 76 76 36 36 Télécopie : 04 76 76 34 52 
      - Cabinet parlementaire 24 Avenue Alsace-Lorraine 38000 Grenoble Téléphone : 04 76 47 67 67 Télécopie : 04 76 56 97 75 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Destot
    place_hemicycle: 543
    autresmandats:
      - Maire de Grenoble, Isère (153298 habitants)
    mails:
      - mdestot@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1116.asp
    profession: Ingénieur
    site_web: http://micheldestot.blogs.com/
    debut_mandat: 20/06/2007
    nom: Michel Destot
    type: depute
  depute_1141:
    place_hemicycle: 602
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1141
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1141.asp
    mails:
      - mdolez@assemblee-nationale.fr
      - contact@marc-dolez.org
    adresses:
      - 57 Rue de Bellain 59500 Douai Téléphone : 03 27 87 60 65 Télécopie : 03 27 87 50 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (17ème)
    groupe:
      - gauche démocrate et républicaine / membre
    site_web: http://www.marc-dolez.net
    profession: Maître de conférences
    debut_mandat: 20/06/2007
    nom_de_famille: Dolez
    nom: Marc Dolez
    type: depute
  depute_1152:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 1152
    extras:
      - conseil de surveillance de l'agence centrale des organismes de sécurité sociale / membre titulaire
      - comité de surveillance du fonds de solidarité vieillesse / membre titulaire
    adresses:
      - 91 Rue d'Angleterre 73000 Chambéry Téléphone : 04 79 68 20 39 Télécopie : 04 79 69 27 09 
      - Mairie BP 348 73103 Aix-les-Bains Téléphone : 04 79 35 07 95 Télécopie : 04 79 35 67 74 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Savoie (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Dord
    place_hemicycle: 264
    autresmandats:
      - Président de la communauté d'agglomération du Lac du Bourget
      - Maire d'Aix-les-Bains, Savoie (25717 habitants)
    mails:
      - dord@blogdord.fr
      - ddord@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1152.asp
    profession: Gérant de société
    site_web: http://www.blogdord.fr
    debut_mandat: 20/06/2007
    nom: Dominique Dord
    type: depute
  depute_1155:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - commission des lois / membre / 
    sexe: H
    id_an: 1155
    extras:
      - conseil d'administration de l'institut national des hautes études de sécurité / membre titulaire
    adresses:
      - BP 138 02005 Laon cedex Téléphone : 03 23 23 24 25 Télécopie : 03 23 23 63 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aisne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: René Dosière
    place_hemicycle: 554
    mails:
      - rdosiere@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1155.asp
    profession: Consultant international
    site_web: http://renedosiere.over-blog.com
    debut_mandat: 20/06/2007
    nom: René Dosière
    type: depute
  depute_1165:
    place_hemicycle: 416
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Vice-président du conseil régional (Ile-de-France)
    sexe: H
    id_an: 1165
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1165.asp
    mails:
      - jdray@assemblee-nationale.fr
    adresses:
      - 130 Avenue Gabriel Péri 91700 Sainte-Geneviève-des-Bois Téléphone : 01 69 25 08 04 Télécopie : 01 69 25 01 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Essonne (10ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Enseignant chercheur
    debut_mandat: 20/06/2007
    nom_de_famille: Dray
    nom: Julien Dray
    type: depute
  depute_1166:
    place_hemicycle: 420
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1166
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1166.asp
    mails:
      - tdreyfus@assemblee-nationale.fr
    adresses:
      - 77  Rue du faubourg Saint-Martin 75010 Paris Téléphone : 01 40 40 40 20 Télécopie : 01 40 40 40 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Avocat au Barreau de Paris
    debut_mandat: 20/06/2007
    nom_de_famille: Dreyfus
    nom: Tony Dreyfus
    type: depute
  depute_1182:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1182
    extras:
      - conférence nationale des services d'incendie et de secours / membre suppléant
    adresses:
      - Mairie 40130 Capbreton Téléphone : 05 58 72 10 09 Télécopie : 05 58 72 25 82 
      - Permanence 1 Rue du Tuc d'Eauze 40100 Dax Téléphone : 05 58 56 09 76 Télécopie : 05 58 56 12 33 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Landes (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Dufau
    place_hemicycle: 362
    autresmandats:
      - Maire de Capbreton, Landes (6678 habitants)
    mails:
      - jpdufau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1182.asp
    profession: Enseignant retraité
    site_web: http://www.jeanpierredufau.org
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Dufau
    type: depute
  depute_1193:
    place_hemicycle: 465
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Premier Vice-président du conseil général (Gard)
    sexe: H
    id_an: 1193
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1193.asp
    mails:
      - dumas.william@wanadoo.fr
      - wdumas@assemblee-nationale.fr
    adresses:
      - 15  Route de Salinelles BP 82012 30252 Sommières cedex Téléphone : 04 66 80 60 60 Télécopie : 04 66 80 60 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gard (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.williamdumas.net
    debut_mandat: 20/06/2007
    nom_de_famille: Dumas
    nom: William Dumas
    type: depute
  depute_1198:
    place_hemicycle: 644
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 1198
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1198.asp
    mails:
      - ejardin-payet.ldumont@orange.fr
      - pleroy.ldumont@orange.fr
      - dumont-laurence@orange.fr
      - ldumont@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 17 Rue Paul Toutain 14000 Caen Téléphone : 02 31 78 15 10 Télécopie : 02 31 72 86 31 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.laurencedumont.net
    profession: Chargée d'études
    debut_mandat: 20/06/2007
    nom_de_famille: Dumont
    nom: Laurence Dumont
    type: depute
  depute_1199:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 1199
    extras:
      - observatoire national du service public de l'électricité et du gaz / membre suppléant
      - conseil de l'immobilier de l'etat / membre titulaire
      - comité local d'information et de suivi du laboratoire souterrain de bure / membre titulaire
      - conseil de surveillance de l'agence française de développement / membre suppléant
    adresses:
      - 7 Rue de la Liberté 55100 Verdun 
      - Permanence 1  Avenue Garibaldi BP 70075 55102 Verdun cedex Téléphone : 03 29 84 85 55 Télécopie : 03 29 84 85 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meuse (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Dumont
    place_hemicycle: 557
    autresmandats:
      - Membre du Conseil municipal de Verdun, Meuse (19621 habitants)
    mails:
      - jldumont@assemblee-nationale.fr
      - Jean-Louis.Dumont@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1199.asp
    profession: Enseignant
    site_web: http://www.jeanlouisdumont.fr
    debut_mandat: 20/06/2007
    nom: Jean-Louis Dumont
    type: depute
  depute_1205:
    place_hemicycle: 114
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Membre du conseil général (Corrèze)
    sexe: H
    id_an: 1205
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1205.asp
    mails:
      - jpdupont@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 3 Rue Saint-Martin 19200 Ussel 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Corrèze (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Docteur vétérinaire
    debut_mandat: 20/06/2007
    nom_de_famille: Dupont
    nom: Jean-Pierre Dupont
    type: depute
  depute_1206:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1206
    adresses:
      - Mairie 60 Rue Charles de Gaulle 91335 Yerres cedex Téléphone : 01 69 49 29 30 Télécopie : 01 69 06 05 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Essonne (8ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    nom_de_famille: Dupont-Aignan
    place_hemicycle: 68
    autresmandats:
      - Maire d'Yerres, Essonne (27457 habitants)
    mails:
      - ndupont@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1206.asp
    profession: Administrateur civil
    site_web: http://www.nicolasdupontaignan.fr
    debut_mandat: 20/06/2007
    nom: Nicolas Dupont-Aignan
    type: depute
  depute_1208:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1208
    adresses:
      - 90 Rue Saint-Martin 11300 Limoux Téléphone : 04 68 31 67 67 Télécopie : 04 68 31 70 70 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville Rue de la Mairie 11300 Limoux Téléphone : 04 68 31 01 16 Télécopie : 04 68 31 85 09 
    circonscription: Aude (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Jean-Paul Dupré
    place_hemicycle: 455
    autresmandats:
      - Maire de Limoux, Aude (9410 habitants)
    mails:
      - jpdupre@assemblee-nationale.fr
      - jp.dupre@ataraxie.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1208.asp
    profession: Cadre bancaire retraité
    site_web: http://www.jean-paul-dupre.fr
    debut_mandat: 20/06/2007
    nom: Jean-Paul Dupré
    type: depute
  depute_1214:
    place_hemicycle: 475
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Maire de Lomme, Nord (27940 habitants)
    sexe: H
    id_an: 1214
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1214.asp
    mails:
      - yvesdurand.lomme@orange.fr
      - ydurand@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 351  Avenue de Dunkerque BP 20415 59464 Lomme cedex Téléphone : 03 20 93 00 59 Télécopie : 03 20 93 97 75 
      - Mairie 59160 Lomme Téléphone : 03 20 22 76 22 Télécopie : 03 20 92 95 88 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (11ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Enseignant
    debut_mandat: 20/06/2007
    nom_de_famille: Durand
    nom: Yves Durand
    type: depute
  depute_1224:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 1224
    adresses:
      - Permanence parlementaire 25  Rue du Bois BP 9 62149 Cambrin Téléphone : 03 21 27 83 29 Télécopie : 03 21 27 91 87 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (11ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Duriez
    place_hemicycle: 511
    autresmandats:
      - Membre du conseil général (Pas-de-Calais)
      - Maire de Cambrin, Pas-de-Calais (957 habitants)
      - Membre de la communauté d'agglomération de l'Artois
    mails:
      - oduriez@assemblee-nationale.fr
      - duriez.odette@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1224.asp
    profession: Comptable
    site_web: http://www.odetteduriez.com
    debut_mandat: 20/06/2007
    nom: Odette Duriez
    type: depute
  depute_1226:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1226
    adresses:
      - Mairie Esplanade Jean-Marie Louvel 14000 Caen Téléphone : 02 31 30 40 50 Télécopie : 02 31 30 45 80 
      - Permanence parlementaire 55 Rue des Jacobins 14000 Caen Téléphone : 02 31 96 49 91 Télécopie : 02 31 77 51 34 
      - Caen la Mer 21 Place de la République 14000 Caen 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Duron
    place_hemicycle: 439
    autresmandats:
      - Président de la communauté d'agglomération de Caen la Mer
      - Maire de Caen, Calvados (114002 habitants)
    mails:
      - philippeduron@orange.fr
      - pduron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1226.asp
    profession: Professeur de lycée agrégé d'histoire
    site_web: http://philippe-duron.fr/blog
    debut_mandat: 20/06/2007
    nom: Philippe Duron
    type: depute
  depute_1243:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 1243
    adresses:
      - 8 Rue Alfred Mézières 54400 Longwy 
      - Hôtel de ville 54750 Trieux 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meurthe-et-Moselle (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Eckert
    place_hemicycle: 648
    autresmandats:
      - Vice-président du conseil régional (Lorraine)
      - Maire de Trieux, Meurthe-et-Moselle (1853 habitants)
    mails:
      - ceckert@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1243.asp
    profession: Professeur
    site_web: http://christianeckert.over-blog.com
    debut_mandat: 20/06/2007
    nom: Christian Eckert
    type: depute
  depute_1252:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 1252
    adresses:
      - Rue de la Paix 40380 Montfort-en-Chalosse Téléphone : 05 58 98 63 70 Télécopie : 05 58 98 57 19 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Landes (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Emmanuelli
    place_hemicycle: 501
    autresmandats:
      - Président du conseil général (Landes)
    mails:
      - hemmanuelli@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1252.asp
    profession: Directeur-adjoint de banque
    site_web: http://www.henriemmanuelli.fr
    debut_mandat: 20/06/2007
    nom: Henri Emmanuelli
    type: depute
  depute_1263:
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Nice, Alpes-Maritimes (342482 habitants)
      - Président de la communauté urbaine Nice - Côte d'Azur
    sexe: H
    id_an: 1263
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1263.asp
    circonscription: Alpes-Maritimes (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Ancien sportif de haut niveau
    debut_mandat: 26/05/2008
    nom_de_famille: Estrosi
    nom: Christian Estrosi
    type: depute
  depute_1268:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1268
    adresses:
      - Mairie Esplanade Tony Larue 76120 Grand-Quevilly Téléphone : 02 35 68 93 00 Télécopie : 02 35 67 27 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Fabius
    place_hemicycle: 515
    autresmandats:
      - Premier adjoint de Grand-Quevilly, Seine-Maritime (26710 habitants)
    mails:
      - lfabius@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1268.asp
    profession: Ancien Maître des requêtes au Conseil d'Etat
    site_web: http://www.laurent-fabius.net
    debut_mandat: 20/06/2007
    nom: Laurent Fabius
    type: depute
  depute_1271:
    place_hemicycle: 512
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Membre du Conseil municipal de Courrières, Pas-de-Calais (10592 habitants)
    sexe: H
    id_an: 1271
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1271.asp
    mails:
      - afacon@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire Place Jean Tailliez 62710 Courrières Téléphone : 03 21 49 11 98 Télécopie : 03 21 49 21 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (14ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur
    debut_mandat: 20/06/2007
    nom_de_famille: Facon
    nom: Albert Facon
    type: depute
  depute_1300:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1300
    adresses:
      - 232 Boulevard Maréchal Leclerc BP 101 84203 Carpentras cedex Téléphone : 04 90 67 10 19 Télécopie : 04 90 63 02 09 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vaucluse (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ferrand
    place_hemicycle: 105
    autresmandats:
      - Membre du conseil général (Vaucluse)
    mails:
      - jmferrand@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1300.asp
    profession: Professeur de lettres
    site_web: http://www.jeanmichelferrand.com
    debut_mandat: 20/06/2007
    nom: Jean-Michel Ferrand
    type: depute
  depute_1304:
    place_hemicycle: 297
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Membre de la Communauté de communes de la Haute Bruche
      - Maire de Wisches, Bas-Rhin (2017 habitants)
    sexe: H
    id_an: 1304
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1304.asp
    mails:
      - alain.ferry2@wanadoo.fr
      - aferry@assemblee-nationale.fr
    adresses:
      - 2 Rue des Ecoles 67130 Wisches Téléphone : 03 88 47 36 45 Télécopie : 03 88 47 39 92 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (6ème)
    groupe:
      - union pour un mouvement populaire / apparenté
    profession: Chef d'entreprise
    debut_mandat: 20/06/2007
    nom_de_famille: Ferry
    nom: Alain Ferry
    type: depute
  depute_1326:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1326
    extras:
      - comité de liaison pour l'accessibilité des transports et du cadre bâti / membre titulaire
    adresses:
      - Permanence parlementaire 1  Rue Émile Péreire 65000 Tarbes Téléphone : 05 62 38 00 42 Télécopie : 05 62 38 09 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hautes-Pyrénées (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Forgues
    place_hemicycle: 474
    autresmandats:
      - Vice-président du conseil régional (Midi-Pyrénées)
    mails:
      - pierre.forgues@laposte.net
      - pforgues@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1326.asp
    profession: Professeur de mathématiques
    debut_mandat: 20/06/2007
    nom: Pierre Forgues
    type: depute
  depute_1327:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 1327
    extras:
      - conférence de la ruralité / membre titulaire
      - conseil supérieur de la participation / membre titulaire
    adresses:
      - 6 Rue des Trois Marchands 36400 La Châtre Téléphone : 02 54 48 02 47 Télécopie : 02 54 48 38 33 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Indre (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Forissier
    place_hemicycle: 344
    autresmandats:
      - Président de la communauté de communes de La-Châtre-et-Sainte-Sévère
      - Maire de La Châtre, Indre (4532 habitants)
    mails:
      - nforissier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1327.asp
    profession: Chef d'entreprise
    debut_mandat: 20/06/2007
    nom: Nicolas Forissier
    type: depute
  depute_1341:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission des finances / membre / 
    sexe: H
    id_an: 1341
    extras:
      - comité des prix de revient des fabrications d'armement / membre titulaire
    adresses:
      - Mairie Place du Général de Gaulle 78990 Élancourt Téléphone : 01 30 66 44 42 Télécopie : 01 30 66 44 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yvelines (11ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Fourgous
    place_hemicycle: 343
    autresmandats:
      - Maire d'Élancourt, Yvelines (28038 habitants)
    mails:
      - jmfourgous@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1341.asp
    profession: Chef d'entreprise
    site_web: http://www.jmfourgous.com
    debut_mandat: 20/06/2007
    nom: Jean-Michel Fourgous
    type: depute
  depute_1353:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 1353
    extras:
      - conseil d'administration de la société nationale de programme "la cinquième" / membre titulaire
    adresses:
      - Hôtel de Ville Place de la Mairie BP 10110 60230 Chambly Cedex Téléphone : 01 39 37 44 13 Télécopie : 01 72 72 96 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Françaix
    place_hemicycle: 457
    autresmandats:
      - Maire de Chambly, Oise (9138 habitants)
    mails:
      - mfrancaix@assemblee-nationale.fr
      - michel.francaix@ville-chambly.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1353.asp
    profession: Consultant en communication
    site_web: http://www.michelfrancaix.fr
    debut_mandat: 20/06/2007
    nom: Michel Françaix
    type: depute
  depute_1355:
    place_hemicycle: 274
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Maire de Puteaux, Hauts-de-Seine (40671 habitants)
    sexe: F
    id_an: 1355
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1355.asp
    mails:
      - jceccaldi@gmail.com
      - jceccaldi@assemblee-nationale.fr
      - joelle.ceccaldi@mairie-puteaux.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie 131 Rue de la République 92801 Puteaux cedex 
    circonscription: Hauts-de-Seine (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Ancien clerc de notaire
    debut_mandat: 20/06/2007
    nom_de_famille: Ceccaldi-Raynaud
    nom: Joëlle Ceccaldi-Raynaud
    type: depute
  depute_1364:
    fonctions:
      - commission des affaires sociales / secrétaire / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 1364
    extras:
      - conseil d'administration de l'établissement d'hospitalisation public de fresnes spécifiquement destine à l'accueil des personnes incarcérées / membre suppléante
    adresses:
      - Hôtel de Ville Rue du 8 Mai 1945 92000 Nanterre Téléphone : 01 70 72 47 24 Télécopie : 01 70 72 47 17 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hauts-de-Seine (4ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Fraysse
    place_hemicycle: 590
    autresmandats:
      - Membre du Conseil municipal de Nanterre, Hauts-de-Seine (84273 habitants)
    mails:
      - jacqueline.fraysse@mairie-nanterre.fr
      - jfraysse@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1364.asp
    profession: Médecin cardiologue
    debut_mandat: 20/06/2007
    nom: Jacqueline Fraysse
    type: depute
  depute_1375:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1375
    extras:
      - comité de l'initiative française pour les récifs coralliens / membre titulaire
    adresses:
      - BP 732 98849 Nouméa cedex 
      - Assemblée de la Province Sud BP L1  Nouméa cedex Téléphone : (687) 25 81 59 Télécopie : (687) 25 81 58 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nouvelle-Calédonie (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Frogier
    place_hemicycle: 277
    autresmandats:
      - Président de l'Assemblée de la province Sud de la Nouvelle Calédonie
    mails:
      - pfrogier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1375.asp
    profession: Administrateur de biens
    debut_mandat: 20/06/2007
    nom: Pierre Frogier
    type: depute
  depute_1379:
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / président / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1379
    extras:
      - commission de vérification des fonds spéciaux (art 154 de la loi de finances pour 2002 / membre titulaire
      - comité des prix de revient des fabrications d'armement / membre titulaire
    adresses:
      - Secrétariat parlementaire Hôtel de ville 18700 Aubigny-sur-Nère Téléphone : 02 48 81 50 91 Télécopie : 02 48 81 50 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Cher (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Fromion
    place_hemicycle: 272
    autresmandats:
      - Vice-président de la Communauté de communes Sauldre et Sologne
      - Maire d'Aubigny-sur-Nère, Cher (5908 habitants)
    mails:
      - yves@fromion.org
      - yfromion@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1379.asp
    profession: Sous-préfet
    site_web: http://www.fromion.org
    debut_mandat: 20/06/2007
    nom: Yves Fromion
    type: depute
  depute_1399:
    place_hemicycle: 3
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire de Saint-Saulve, Nord (11027 habitants)
    sexe: F
    id_an: 1399
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1399.asp
    circonscription: Nord (21ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Pharmacienne retraitée
    debut_mandat: 20/07/2007
    nom_de_famille: Gallez
    nom: Cécile Gallez
    type: depute
  depute_1418:
    place_hemicycle: 148
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 1418
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1418.asp
    mails:
      - garrigue.daniel.depute@wanadoo.fr
      - dgarrigue@assemblee-nationale.fr
    adresses:
      - Permanence 2 Rue des 2 conils 24100 Bergerac Téléphone : 05 53 27 65 35 Télécopie : 05 53 58 22 31 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Dordogne (2ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    site_web: http://www.danielgarrigue.com
    profession: Administrateur à l'Assemblée nationale
    debut_mandat: 20/06/2007
    nom_de_famille: Garrigue
    nom: Daniel Garrigue
    type: depute
  depute_1432:
    place_hemicycle: 261
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1432
    extras:
      - haut comité pour la transparence et l'information sur la sécurité nucléaire / membre titulaire
      - observatoire national du service public de l'électricité et du gaz / membre titulaire
      - haut conseil des biotechnologies / membre titulaire
      - conseil supérieur de l'aviation marchande / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1432.asp
    mails:
      - claude.gatignol.permanence@wanadoo.fr
      - cgatignol@assemblee-nationale.fr
    adresses:
      - 2 Rue des Résistants 50700 Valognes Téléphone : 02 33 95 15 00 Télécopie : 02 33 95 13 57 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Manche (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Docteur vétérinaire
    debut_mandat: 20/06/2007
    nom_de_famille: Gatignol
    nom: Claude Gatignol
    type: depute
  depute_1433:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / vice-président / 
    sexe: H
    id_an: 1433
    extras:
      - commission nationale de présélection des pôles d'excellence rurale / membre titulaire
      - observatoire national du service public de l'électricité et du gaz / membre suppléant
    adresses:
      - 12 Bis Rue de Brest 22100 Dinan Téléphone : 02 96 39 09 50 Télécopie : 02 96 39 19 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 04 06 Télécopie : 01 40 63 04 86 
    circonscription: Côtes-d'Armor (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Gaubert
    place_hemicycle: 471
    mails:
      - jgaubert@assemblee-nationale.fr
      - jean-gaubert@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1433.asp
    profession: Agriculteur-éleveur
    site_web: http://jeangaubert.typepad.com
    debut_mandat: 20/06/2007
    nom: Jean Gaubert
    type: depute
  depute_1445:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1445
    extras:
      - conseil supérieur des archives / membre titulaire
    adresses:
      - 5 Place Ferdinand Million 73200 Albertville Téléphone : 04 79 32 03 68 Télécopie : 04 79 37 82 74 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Savoie (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gaymard
    place_hemicycle: 170
    autresmandats:
      - Président du conseil général (Savoie)
    mails:
      - hgaymard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1445.asp
    profession: Administrateur civil
    debut_mandat: 20/06/2007
    nom: Hervé Gaymard
    type: depute
  depute_1452:
    fonctions:
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
      - commission des affaires sociales / vice-présidente / 
    sexe: F
    id_an: 1452
    extras:
      - conseil de modération et de prévention / membre titulaire
    adresses:
      - 70 Rue des Trois Visages 62000 Arras Téléphone : 03 21 73 51 66 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Génisson
    place_hemicycle: 496
    autresmandats:
      - Vice-présidente du conseil régional (Nord-Pas-de-Calais)
    mails:
      - cgenisson@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1452.asp
    profession: Praticien hospitalier
    site_web: http://www.catherine-genisson.fr
    debut_mandat: 20/06/2007
    nom: Catherine Génisson
    type: depute
  depute_1459:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1459
    extras:
      - conseil d'administration de l'établissement public national d'aménagement et de restructuration des espaces commerciaux et artisanaux / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 103 Avenue Foch 59700 Marcq-en-Baroeul Téléphone : 08 10 45 45 45 Télécopie : 03 20 45 45 37 
    circonscription: Nord (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gérard
    place_hemicycle: 324
    autresmandats:
      - Maire de Marcq-en-Baroeul, Nord (37174 habitants)
    mails:
      - bgerard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1459.asp
    profession: Avocat
    debut_mandat: 20/06/2007
    nom: Bernard Gérard
    type: depute
  depute_1463:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1463
    adresses:
      - Permanence parlementaire 27 Rue Francis de Préssensé 69190 Saint-Fons Téléphone : 04 78 67 16 99 Télécopie : 04 78 67 16 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville 5  Avenue Marcel Houel BP 24 69631 Vénissieux cedex Téléphone : 04 72 21 44 68 Télécopie : 04 72 21 45 02 
    circonscription: Rhône (14ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Gerin
    place_hemicycle: 576
    autresmandats:
      - Maire de Vénissieux, Rhône (56061 habitants)
    mails:
      - andregerin@orange.fr
      - agerin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1463.asp
    profession: Dessinateur industriel
    site_web: http://www.andregerin.com
    debut_mandat: 20/06/2007
    nom: André Gerin
    type: depute
  depute_1466:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / secrétaire / 
      - délégation chargée de la communication et de la presse / membre / 
      - assemblée nationale / secrétaire / 01/10/2008
    sexe: H
    id_an: 1466
    extras:
      - conseil d'orientation pour la prévention des risques naturels majeurs / membre titulaire
    adresses:
      - 32 Rue Jules Lardière 80800 Corbie Téléphone : 03 22 96 07 68 Télécopie : 03 22 96 07 69 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Somme (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gest
    place_hemicycle: 260
    mails:
      - agest@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1466.asp
    profession: Consultant
    site_web: http://www.alaingest.info
    debut_mandat: 20/06/2007
    nom: Alain Gest
    type: depute
  depute_1477:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 1477
    extras:
      - comité d'enquête sur le coût et le rendement des services publics / membre titulaire
      - conférence nationale des services d'incendie et de secours / membre titulaire
    adresses:
      - Permanence parlementaire 60  Allée Frédéric Mistral Boulouris 83700 Saint-Raphaël 
      - Hôtel de Ville BP 80160 83701 Saint-Raphaël cedex Téléphone : 04 94 82 15 17 Télécopie : 04 94 19 19 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Var (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ginesta
    place_hemicycle: 313
    autresmandats:
      - Président de la communauté d'agglomération de Fréjus-Saint-Raphaël
      - Maire de Saint-Raphaël, Var (30664 habitants)
    mails:
      - gginesta@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1477.asp
    profession: Ingénieur ETP
    debut_mandat: 20/06/2007
    nom: Georges Ginesta
    type: depute
  depute_1483:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1483
    extras:
      - conseil d'administration des parcs nationaux de france / membre titulaire
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 14 Rue Jean Aicard 83400 Hyères Téléphone : 04 94 65 64 49 Télécopie : 04 94 65 73 42 
    circonscription: Var (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Giran
    place_hemicycle: 102
    autresmandats:
      - Membre du Conseil municipal de Hyères, Var (51417 habitants)
    mails:
      - jeanpierre.giran@wanadoo.fr
      - jpgiran@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1483.asp
    profession: Professeur d'Université
    site_web: http://www.giran.fr
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Giran
    type: depute
  depute_1496:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1496
    adresses:
      - Permanence 170 Place de la Libération 65700 Maubourguet Téléphone : 05 62 96 99 27 Télécopie : 05 62 96 39 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 94 19 
    circonscription: Hautes-Pyrénées (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Glavany
    place_hemicycle: 495
    autresmandats:
      - Membre du Conseil municipal de Tarbes, Hautes-Pyrénées (46275 habitants)
    mails:
      - glavany.jean@wanadoo.fr
      - jglavany@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1496.asp
    profession: Préfet
    site_web: http://www.jean-glavany.net
    debut_mandat: 20/06/2007
    nom: Jean Glavany
    type: depute
  depute_1498:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / vice-président / 
      - commission des lois / membre / 
    sexe: H
    id_an: 1498
    extras:
      - commission nationale de l'admission exceptionnelle au séjour / membre titulaire
    adresses:
      - Mairie de Paris 9 Place de l'Hôtel de Ville 75196 Paris RP Téléphone : 01 42 76 65 46 Télécopie : 01 42 76 46 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (14ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Goasguen
    place_hemicycle: 172
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Maire d'arrondissement de Paris (16ème Arrondissement), Paris (160007 habitants)
      - Conseiller de Paris
    mails:
      - cgoasguen@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1498.asp
    profession: Avocat à la Cour d'appel de Paris
    site_web: http://www.claudegoasguen.typepad.com
    debut_mandat: 20/06/2007
    nom: Claude Goasguen
    type: depute
  depute_1514:
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1514
    extras:
      - conseil national des transports / membre titulaire
    adresses:
      - Permanence parlementaire 40 Ter Rue Saint Eloi 60400 NOYON Téléphone : 03 44 09 12 19 Télécopie : 03 44 09 12 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gonnot
    place_hemicycle: 258
    autresmandats:
      - Membre du Conseil municipal de Noyon, Oise (14471 habitants)
    mails:
      - fmgonnot@assemblee-nationale.fr
      - gonnot2007@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1514.asp
    profession: Conseil en entreprises
    site_web: http://gonnot.over-blog.com
    debut_mandat: 20/06/2007
    nom: François-Michel Gonnot
    type: depute
  depute_1515:
    fonctions:
      - commission des affaires étrangères / membre / 
      - mission d'évaluation de la loi n°2005-370 du 22 avril 2005 relative aux droits des malades et à la fin de vie / membre / 
      - mission d'information commune sur les exonérations sociales / membre / 
    sexe: H
    id_an: 1515
    extras:
      - conseil d'orientation pour l'emploi / membre titulaire
    adresses:
      - 9 Rue Saint-Jacques 58200 Cosne-sur-Loire Téléphone : 03 86 26 91 99 Télécopie : 03 86 26 89 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nièvre (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Gorce
    place_hemicycle: 423
    autresmandats:
      - Maire de la Charité-sur-Loire, Nièvre (5460 habitants)
    mails:
      - ggorce@assemblee-nationale.fr
      - GORCE.GAETAN@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1515.asp
    profession: Administrateur civil
    site_web: http://gorce.typepad.fr/blog/
    debut_mandat: 20/06/2007
    nom: Gaëtan Gorce
    type: depute
  depute_1521:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 1521
    extras:
      - commission nationale des compétences et des talents / membre titulaire
      - conseil d'orientation de l'observatoire national de la délinquance / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 00 
      - Mairie du 15ème Rue Peclet 75015 Paris Téléphone : 01 55 76 75 00 Télécopie : 01 55 76 75 18 
    circonscription: Paris (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Goujon
    place_hemicycle: 232
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Maire d'arrondissement de Paris (15ème Arrondissement), Paris (225410 habitants)
      - Conseiller de Paris
    mails:
      - pgoujon@assemblee-nationale.fr
      - philippegoujon@hotmail.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1521.asp
    profession: Cadre
    debut_mandat: 20/06/2007
    nom: Philippe Goujon
    type: depute
  depute_1522:
    place_hemicycle: 255
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Maire de Vannes, Morbihan (51759 habitants)
      - Président de la communauté d'agglomération du Pays de Vannes
    sexe: H
    id_an: 1522
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1522.asp
    mails:
      - fgoulard@assemblee-nationale.fr
    adresses:
      - Permanence 2 Rue de la Boucherie 56000 VANNES Téléphone : 02 97 47 05 10 Télécopie : 02 97 47 80 13 
      - Hôtel de ville Place Maurice Marchais 56000 Vannes Téléphone : 02 97 01 60 10 Télécopie : 02 97 01 60 11 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Morbihan (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.fgoulard.fr
    debut_mandat: 20/06/2007
    nom_de_famille: Goulard
    nom: François Goulard
    type: depute
  depute_1548:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 1548
    extras:
      - conseil d'orientation des retraites / membre titulaire
      - comité national des retraités et des personnes âgées / membre suppléant
      - conseil national de la formation professionnelle tout au long de la vie / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 39 Rue Lamarck 80000 Amiens Téléphone : 03 22 97 35 53 Télécopie : 03 22 97 39 04 
      - 16 Rue Gaudissart 80000 Amiens Téléphone : 03 22 91 78 44 Télécopie : 03 22 92 87 24 
    circonscription: Somme (1ère)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Gremetz
    place_hemicycle: 595
    autresmandats:
      - Membre du conseil régional (Picardie)
    mails:
      - contact@maxime-gremetz.fr
      - mgremetz@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1548.asp
    profession: Métallurgiste
    site_web: http://www.maxime-gremetz.fr
    debut_mandat: 20/06/2007
    nom: Maxime Gremetz
    type: depute
  depute_1549:
    place_hemicycle: 311
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Maire de Bayonne, Pyrénées-Atlantiques (40016 habitants)
    sexe: H
    id_an: 1549
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1549.asp
    mails:
      - jeangrenetdepute@gmail.com
      - jgrenet@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 15 Avenue Foch 64100 Bayonne Téléphone : 05 59 46 24 50 Télécopie : 05 59 46 24 54 
    circonscription: Pyrénées-Atlantiques (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chirurgien retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Grenet
    nom: Jean Grenet
    type: depute
  depute_1562:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / secrétaire / 
    sexe: H
    id_an: 1562
    adresses:
      - Permanence parlementaire 57140 Woippy Téléphone : 03 87 30 44 15 Télécopie : 03 87 30 74 87 
      - Mairie 57140 Woippy Téléphone : 03 87 34 63 42 Télécopie : 03 87 34 63 33 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Moselle (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Grosdidier
    place_hemicycle: 215
    autresmandats:
      - Maire de Woippy, Moselle (13755 habitants)
    mails:
      - fgrosdidier@assemblee-nationale.fr
      - woippy.grosdidier@wanadoo.fr
      - permanence.francoisgrosdidier@voila.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1562.asp
    profession: Fonctionnaire territorial
    site_web: http://www.fgrosdidier.fr
    debut_mandat: 20/06/2007
    nom: François Grosdidier
    type: depute
  depute_1568:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1568
    extras:
      - conseil national du littoral / membre titulaire
      - conseil de surveillance de l'agence française de développement / membre suppléant
    adresses:
      - Hôtel de Ville BP 30386 85108 Les Sables-d'Olonne Téléphone : 02 51 23 16 02 
      - 40 Rue de Bel Air 85100 Les Sables d'Olonne Téléphone : 08 79 57 04 31 Télécopie : 02 51 21 58 87 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vendée (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Guédon
    place_hemicycle: 213
    autresmandats:
      - Maire des Sables-d'Olonne, Vendée (15532 habitants)
      - Président de la communauté de communes des Olonnes
    mails:
      - lguedon@assemblee-nationale.fr
      - louis.guedon885@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1568.asp
    profession: Docteur en  pharmacie, biologiste
    debut_mandat: 20/06/2007
    nom: Louis Guédon
    type: depute
  depute_1574:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1574
    extras:
      - conseil national du littoral / membre titulaire
    adresses:
      - Permanence 7 Place de la Mairie 06500 Menton Téléphone : 09 54 10 86 13 Télécopie : 04 93 41 38 06 
      - Hôtel de Ville 17 Rue de la République 06500 Menton 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-Maritimes (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Guibal
    place_hemicycle: 187
    autresmandats:
      - Maire de Menton, Alpes-Maritimes (28862 habitants)
    mails:
      - jcguibal@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1574.asp
    profession: Ancien dirigeant d'organisations professionnelles
    debut_mandat: 20/06/2007
    nom: Jean-Claude Guibal
    type: depute
  depute_1579:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: F
    id_an: 1579
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 93 20 Télécopie : 01 40 63 93 36 
      - BP 47 93141 Bondy cedex Téléphone : 01 48 50 04 67 Télécopie : 01 48 49 66 72 
    circonscription: Seine-Saint-Denis (9ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Guigou
    place_hemicycle: 412
    autresmandats:
      - Adjointe au Maire de Noisy-le-Sec, Seine-Saint-Denis (37312 habitants)
    mails:
      - eguigou@assemblee-nationale.fr
      - guigou.e@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1579.asp
    profession: Administrateur civil du ministère des finances
    site_web: http://elisabethguigou.hautetfort.com
    debut_mandat: 20/06/2007
    nom: Élisabeth Guigou
    type: depute
  depute_1585:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1585
    adresses:
      - 2 Bis Avenue de l'Europe 92310 Sèvres Téléphone : 01 45 34 09 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hauts-de-Seine (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Guillet
    place_hemicycle: 165
    autresmandats:
      - Premier vice-président de la communauté d'agglomération Arc de Seine
      - Maire de Chaville, Hauts-de-Seine (17939 habitants)
    mails:
      - jjguillet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1585.asp
    profession: Chef d'entreprise retraité
    site_web: http://www.jjguillet.org
    debut_mandat: 20/06/2007
    nom: Jean-Jacques Guillet
    type: depute
  depute_1592:
    place_hemicycle: 446
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / coprésident / 
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission des finances / membre / 
    autresmandats:
      - Président de la communauté de communes de Lacq
      - Maire de Mourenx, Pyrénées-Atlantiques (7537 habitants)
    sexe: H
    id_an: 1592
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1592.asp
    mails:
      - dhabib.orthez@wanadoo.fr
      - dhabib@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 51 Rue Saint-Gilles 64300 Orthez Téléphone : 05 59 67 20 07 Télécopie : 05 59 67 20 02 
      - Mairie Place François Mitterrand 64150 Mourenx Téléphone : 05 59 60 07 23 Télécopie : 05 59 60 07 90 
      - Hôtel de la Communauté de communes Rond-Point des Chênes 64150 Mourenx Téléphone : 05 59 60 03 46  Télécopie : 05 59 60 95 43 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Atlantiques (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre
    debut_mandat: 20/06/2007
    nom_de_famille: Habib
    nom: David Habib
    type: depute
  depute_1604:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1604
    extras:
      - conseil d'administration de l'agence nationale pour la cohésion sociale et l'égalité des chances / membre titulaire
      - commission nationale chargée de l'examen du respect des obligations de réalisation de logements sociaux / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 67 95 Télécopie : 01 40 63 56 91 
      - Permanence parlementaire 33 Boulevard Louis Terrier 28100 Dreux Téléphone : 02 37 50 10 41 Télécopie : 02 37 50 11 22 
      - Mairie 2 Rue de Châteaudun BP 129 28103 Dreux cedex Téléphone : 02 37 38 84 45 Télécopie : 02 37 38 84 05 
    circonscription: Eure-et-Loir (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Hamel
    place_hemicycle: 251
    autresmandats:
      - Maire de Dreux, Eure-et-Loir (31898 habitants)
      - Président Communauté d'Agglomération du Drouais
    mails:
      - g.hamel@ville-dreux.fr
      - ghamel@assemblee-nationale.fr
      - permanence.ghamel@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1604.asp
    profession: Chef d'entreprise du bâtiment
    debut_mandat: 20/06/2007
    nom: Gérard Hamel
    type: depute
  depute_1630:
    fonctions:
      - commission des affaires culturelles et de l'éducation / vice-président / 
      - commission des affaires européennes / vice-président / 
    sexe: H
    id_an: 1630
    extras:
      - conseil d'administration de l'agence pour l'enseignement français à l'étranger / membre suppléant
      - comité de suivi de la mise en oeuvre des dispositions relatives au cinéma et autres arts et industries de l'image animée / membre titulaire
      - conseil d'administration de la société en charge de l'audiovisuel extérieur de la france / membre titulaire
      - conseil d'administration du centre national d'art et de culture georges pompidou / membre titulaire
      - conseil d'administration de l'hôpital national de saint-maurice / membre titulaire
    adresses:
      - Hôtel de Ville 118 Avenue du Général de Gaulle 94700 Maisons-Alfort Téléphone : 01 43 96 77 23 Télécopie : 01 43 96 96 38 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Herbillon
    place_hemicycle: 259
    autresmandats:
      - Maire de Maisons-Alfort, Val-de-Marne (54000 habitants)
    mails:
      - mherbillon@assemblee-nationale.fr
      - michel.herbillon@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1630.asp
    profession: Cadre
    site_web: http://www.maisons-alfort.fr
    debut_mandat: 20/06/2007
    nom: Michel Herbillon
    type: depute
  depute_1654:
    place_hemicycle: 509
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Président du conseil général (Corrèze)
    sexe: H
    id_an: 1654
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1654.asp
    mails:
      - fhollande@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 36 Avenue Victor Hugo 19000 Tulle Téléphone : 05 55 20 48 48 Télécopie : 05 55 20 38 38 
    circonscription: Corrèze (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Conseiller référendaire à la Cour des comptes
    debut_mandat: 20/06/2007
    nom_de_famille: Hollande
    nom: François Hollande
    type: depute
  depute_1658:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: F
    id_an: 1658
    adresses:
      - BP 97 59850 Nieppe Téléphone : 03 20 57 31 86 Télécopie : 03 20 57 36 92 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (15ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Hostalier
    place_hemicycle: 64
    autresmandats:
      - Membre du conseil régional (Nord-Pas-de-Calais)
    mails:
      - fhostalier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1658.asp
    profession: Inspecteur général de l'Education nationale
    site_web: http://www.francoisehostalier.fr
    debut_mandat: 20/06/2007
    nom: Françoise Hostalier
    type: depute
  depute_1661:
    place_hemicycle: 337
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Pontoise, Val-d'Oise (27477 habitants)
    sexe: H
    id_an: 1661
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1661.asp
    mails:
      - phouillon@assemblee-nationale.fr
    adresses:
      - Permanence 11 Place de l'Hôtel de Ville 95300 Pontoise Téléphone : 01 30 38 55 89 Télécopie : 01 30 73 11 13 
      - Mairie 2 Rue Victor Hugo 95300 Pontoise Téléphone : 01 34 43 34 43 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Avocat, ancien Bâtonnier de l'Ordre
    debut_mandat: 20/06/2007
    nom_de_famille: Houillon
    nom: Philippe Houillon
    type: depute
  depute_1677:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission des lois / membre / 
    sexe: H
    id_an: 1677
    extras:
      - commission d'accès aux documents administratifs / membre suppléant
      - commission de suivi du mémorandum d'accord signe le 26 novembre 1996 entre la france et la fédération de russie / membre titulaire
      - conseil supérieur de l' administration pénitentiaire / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 11 Place de la Motte 44100 Châteaubriant Téléphone : 02 40 81 45 46 Télécopie : 02 40 81 45 16 
    circonscription: Loire-Atlantique (6ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Hunault
    place_hemicycle: 378
    autresmandats:
      - Membre du conseil régional (Pays de la Loire)
    mails:
      - michel.hunault-depute@wanadoo.fr
      - mhunault@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1677.asp
    profession: Avocat
    site_web: http://www.michel-hunault.com
    debut_mandat: 20/06/2007
    nom: Michel Hunault
    type: depute
  depute_1686:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 1686
    extras:
      - commission centrale de classement des débits de tabac / membre titulaire
      - conseil d'administration de l'office franco-allemand pour la jeunesse / membre suppléant
    adresses:
      - 5 Place Jean Jaurès 31800 Saint-Gaudens Téléphone : 05 62 00 80 80 Télécopie : 05 61 95 99 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Idiart
    place_hemicycle: 541
    autresmandats:
      - Membre du conseil général (Haute-Garonne)
    mails:
      - jean-louis.idiart@wanadoo.fr
      - jlidiart@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1686.asp
    profession: Contrôleur des impôts
    debut_mandat: 20/06/2007
    nom: Jean-Louis Idiart
    type: depute
  depute_1689:
    place_hemicycle: 532
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du conseil régional (Midi-Pyrénées)
    sexe: F
    id_an: 1689
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1689.asp
    mails:
      - fimbert@assemblee-nationale.fr
      - imbert.francoise@wanadoo.fr
    adresses:
      - 17 Allée des Mauges BP 122 31772 Colomiers cedex Téléphone : 05 61 78 61 85 Télécopie : 05 61 78 61 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Ancien chef de cabinet du maire de Colomiers
    debut_mandat: 20/06/2007
    nom_de_famille: Imbert
    nom: Françoise Imbert
    type: depute
  depute_1695:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission du développement durable et de l'aménagement du territoire / président / 
    sexe: H
    id_an: 1695
    adresses:
      - Hôtel de Ville 77160 Provins Téléphone : 01 64 60 38 33 Télécopie : 01 64 00 61 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-et-Marne (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Jacob
    place_hemicycle: 90
    autresmandats:
      - Maire de Provins, Seine-et-Marne (11667 habitants)
      - Président de la communauté de communes du Provinois
    mails:
      - cjacob@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1695.asp
    profession: Agriculteur
    site_web: http://www.christianjacob.fr
    debut_mandat: 20/06/2007
    nom: Christian Jacob
    type: depute
  depute_1699:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 1699
    extras:
      - commission nationale de concertation sur les risques miniers / membre titulaire
      - conseil de surveillance de la caisse nationale d'assurance vieillesse des travailleurs salariés / membre titulaire
      - conseil d'orientation des retraites / membre titulaire
    adresses:
      - Permanence parlementaire 25  Rue du Cambout 57000 Metz Téléphone : 03 87 36 48 28 Télécopie : 03 87 36 11 91 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Moselle (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Jacquat
    place_hemicycle: 135
    autresmandats:
      - Membre du Conseil municipal de Metz, Moselle (123776 habitants)
      - Membre de la communauté d'agglomération de Metz Métropole (CA2M)
    mails:
      - djacquat@wanadoo.fr
      - djacquat@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1699.asp
    profession: Médecin O.R.L.
    site_web: http://www.denisjacquat.fr
    debut_mandat: 20/06/2007
    nom: Denis Jacquat
    type: depute
  depute_1710:
    place_hemicycle: 442
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Membre du Conseil municipal de Bruay-la-Buissière, Pas-de-Calais (23997 habitants)
    sexe: H
    id_an: 1710
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1710.asp
    mails:
      - sjanquin@assemblee-nationale.fr
    adresses:
      - 300 Rue de Vaudricourt 62700 Bruay la Buissière Téléphone : 03 91 80 44 95 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (10ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur certifié de sciences économiques et sociales, enseignement secondaire
    debut_mandat: 20/06/2007
    nom_de_famille: Janquin
    nom: Serge Janquin
    type: depute
  depute_1712:
    fonctions:
      - commission des affaires culturelles et de l'éducation / vice-président / 
      - mission d'évaluation de la loi n°2005-370 du 22 avril 2005 relative aux droits des malades et à la fin de vie / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 1712
    adresses:
      - 103 Ter Rue Victor Hugo 80440 Boves Téléphone : 03 22 09 31 31 Télécopie : 03 22 09 31 31 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Somme (2ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Olivier Jardé
    place_hemicycle: 400
    autresmandats:
      - Membre du conseil général (Somme)
    mails:
      - ojarde@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1712.asp
    profession: Professeur de chirurgie, professeur de droit de la santé
    site_web: http://www.olivierjarde.info
    debut_mandat: 20/06/2007
    nom: Olivier Jardé
    type: depute
  depute_1746:
    place_hemicycle: 16
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1746
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1746.asp
    mails:
      - djulia@assemblee-nationale.fr
      - contact@didier-julia.org
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 67 73 Télécopie : 01 40 63 53 45 
      - Permanence 202 Rue Grande 77300 Fontainebleau Téléphone : 01 64 22 46 30 Télécopie : 01 60 72 33 97 
    circonscription: Seine-et-Marne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Professeur d'Université
    debut_mandat: 20/06/2007
    nom_de_famille: Julia
    nom: Didier Julia
    type: depute
  depute_1748:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1748
    extras:
      - conseil national des transports / membre suppléant
    adresses:
      - 40 Avenue des Vosges 67000 Strasbourg Téléphone : 03 88 24 73 00 Télécopie : 03 88 24 73 03 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Jung
    place_hemicycle: 472
    autresmandats:
      - Membre du conseil général (Bas-Rhin)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1748.asp
    mails:
      - contact@armandjung-depute.fr
    site_web: http://www.armandjung-depute.fr 
    profession: Fonctionnaire territorial
    debut_mandat: 20/06/2007
    nom: Armand Jung
    type: depute
  depute_1761:
    fonctions:
      - commission des affaires culturelles et de l'éducation / vice-président / 
    sexe: H
    id_an: 1761
    extras:
      - conseil d'administration de la société france télévision / membre titulaire
      - conseil d'administration de la fondation du patrimoine / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 14 Rue des Cordeliers 13300 Salon-de-Provence Téléphone : 04 90 56 12 25 Télécopie : 04 90 56 39 98 
    circonscription: Bouches-du-Rhône (11ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Kert
    place_hemicycle: 183
    mails:
      - ckert@assemblee-nationale.fr
      - ckert.cabparlementaire@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1761.asp
    profession: Cadre administratif
    site_web: http://www.christiankert.over-blog.fr
    debut_mandat: 20/06/2007
    nom: Christian Kert
    type: depute
  depute_1770:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1770
    extras:
      - commission de surveillance et de contrôle des publications destinées à l'enfance et à l'adolescence / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville 92401 Courbevoie cedex Téléphone : 01 43 34 70 33 Télécopie : 01 43 34 70 38 
    circonscription: Hauts-de-Seine (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Kossowski
    place_hemicycle: 91
    autresmandats:
      - Maire de Courbevoie, Hauts-de-Seine (68942 habitants)
    mails:
      - jkossowski@assemblee-nationale.fr
      - jakossowski@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1770.asp
    profession: Dirigeant d'entreprise
    site_web: http://quinquasplus.com
    debut_mandat: 20/06/2007
    nom: Jacques Kossowski
    type: depute
  depute_1774:
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - commission des affaires étrangères / secrétaire / 
      - assemblée nationale / secrétaire / 01/10/2008
    sexe: H
    id_an: 1774
    adresses:
      - Centre adminis.- Les Grands Bureaux 45 Rue Edouard Vaillant BP 49 62801 Liévin Téléphone : 03 21 44 89 34 Télécopie : 03 21 44 89 35 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (12ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Kucheida
    place_hemicycle: 507
    autresmandats:
      - Maire de Liévin, Pas-de-Calais (33429 habitants)
    mails:
      - jpkucheida@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1774.asp
    profession: Professeur certifié
    site_web: http://www.jpkucheida.fr/
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Kucheida
    type: depute
  depute_1778:
    place_hemicycle: 13
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Membre du Conseil municipal de Valence, Drôme (64329 habitants)
    sexe: H
    id_an: 1778
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1778.asp
    mails:
      - patrick.labaune@orange.fr
      - plabaune@assemblee-nationale.fr
    adresses:
      - 158 Avenue Victor Hugo Immeuble le Saint Joseph 26000 Valence Téléphone : 09 64 23 81 69 Télécopie : 04 75 42 76 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Drôme (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Enseignant
    debut_mandat: 20/06/2007
    nom_de_famille: Labaune
    nom: Patrick Labaune
    type: depute
  depute_1789:
    place_hemicycle: 531
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Membre de la communauté urbaine de Bordeaux
      - Maire de Floirac, Gironde (16164 habitants)
    sexe: F
    id_an: 1789
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1789.asp
    mails:
      - clacuey@assemblee-nationale.fr
      - clacuey@wanadoo.fr
    adresses:
      - Hôtel de Ville 6 Avenue Pasteur 33270 Floirac Téléphone : 05 57 80 87 44 Télécopie : 05 56 86 77 41 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre comptable
    debut_mandat: 20/06/2007
    nom_de_famille: Lacuey
    nom: Conchita Lacuey
    type: depute
  depute_1790:
    fonctions:
      - commission des affaires européennes / membre / 
      - assemblée nationale / vice-président / 27/06/2007
      - commission des finances / membre / 
      - délégation chargée des activités internationales / président / 
    sexe: H
    id_an: 1790
    extras:
      - comité des finances locales / membre suppléant
      - commission nationale de présélection des pôles d'excellence rurale / membre titulaire
      - conseil de surveillance du fonds de réserve pour les retraites / membre titulaire
    adresses:
      - Cabinet parlementaire Mairie 49240 Avrillé Téléphone : 02 41 37 41 09 Télécopie : 02 41 69 66 41 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 51 78 Télécopie : 01 40 63 97 87 
    circonscription: Maine-et-Loire (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Laffineur
    place_hemicycle: 254
    autresmandats:
      - Maire d'Avrillé, Maine-et-Loire (12991 habitants)
    mails:
      - contact@marclaffineur.org
      - mlaffineur@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1790.asp
    profession: Médecin anesthésiste-réanimateur
    site_web: http://www.marclaffineur.org
    debut_mandat: 20/06/2007
    nom: Marc Laffineur
    type: depute
  depute_1809:
    place_hemicycle: 548
    fonctions:
      - commission des affaires européennes / vice-président / 
      - commission des lois / membre / 
    sexe: H
    id_an: 1809
    extras:
      - commission de surveillance et de contrôle des publications destinées à l'enfance et à l'adolescence / membre suppléant
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1809.asp
    mails:
      - jlambert@assemblee-nationale.fr
    adresses:
      - Le Bourg 16230 Juillé Téléphone : 05 45 39 00 09 Télécopie : 05 45 39 91 74 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Charente (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre de l'industrie
    debut_mandat: 20/06/2007
    nom_de_famille: Lambert
    nom: Jérôme Lambert
    type: depute
  depute_1816:
    place_hemicycle: 497
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Palaiseau, Essonne (28965 habitants)
      - Président de la communauté d'agglomération du Plateau de Saclay
    sexe: H
    id_an: 1816
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1816.asp
    mails:
      - flamy@assemblee-nationale.fr
      - contact@francois-lamy.org
    adresses:
      - Permanence 91 Rue de Paris 91120 Palaiseau Téléphone : 01 60 11 25 77 Télécopie : 01 69 30 71 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 63 Télécopie : 01 40 63 68 50 
    circonscription: Essonne (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Instituteur
    debut_mandat: 20/06/2007
    nom_de_famille: Lamy
    nom: François Lamy
    type: depute
  depute_1821:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1821
    adresses:
      - Permanence parlementaire 74 Rue du Chemin Vert 62200 Boulogne-sur-Mer Téléphone : 03 21 30 91 21 Télécopie : 03 21 30 91 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lang
    place_hemicycle: 419
    autresmandats:
      - Vice-président du conseil régional (Nord-Pas-de-Calais)
    mails:
      - jacklang62@wanadoo.fr
      - jlang@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1821.asp
    profession: Professeur agrégé de droit public
    site_web: http://www.jacklang.org
    debut_mandat: 20/06/2007
    nom: Jack Lang
    type: depute
  depute_1822:
    place_hemicycle: 9
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Maire de Freyming-Merlebach, Moselle (14508 habitants)
      - Président de la Communauté de communes de Freyming-Merlebach
    sexe: H
    id_an: 1822
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1822.asp
    mails:
      - pierrelang@wanadoo.fr
      - plang@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville 42 Rue Nicolas Colson BP 40062 57803 Freyming-Merlebach cedex Téléphone : 03 87 90 59 33 Télécopie : 03 87 90 59 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Moselle (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Biologiste, directeur d'un laboratoire d'analyses médicales
    debut_mandat: 20/06/2007
    nom_de_famille: Lang
    nom: Pierre Lang
    type: depute
  depute_1835:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1835
    extras:
      - conseil de l'agence d'évaluation de la recherche et de l'enseignement supérieur / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 8 Rue Neuve 91190 Gif-sur-Yvette Téléphone : 01 69 28 00 00 Télécopie : 01 69 28 50 07 
    circonscription: Essonne (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lasbordes
    place_hemicycle: 333
    autresmandats:
      - Membre du conseil régional (Ile-de-France)
    mails:
      - p.lasbordes@wanadoo.fr
      - plasbordes@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1835.asp
    profession: Directeur commercial
    site_web: http://www.lasbordes.fr
    debut_mandat: 20/06/2007
    nom: Pierre Lasbordes
    type: depute
  depute_1838:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1838
    extras:
      - conseil national de sécurité civile / membre suppléant
      - commission nationale du débat public  / membre titulaire
    adresses:
      - Permanence 2  Rue Saint-Grat 64400 Oloron-Sainte-Marie Téléphone : 05 59 39 67 83 Télécopie : 05 59 39 06 95 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Atlantiques (4ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    nom_de_famille: Lassalle
    place_hemicycle: 71
    autresmandats:
      - Maire de Lourdios-Ichère, Pyrénées-Atlantiques (150 habitants)
      - Membre du conseil général (Pyrénées-Atlantiques)
    mails:
      - jlassalle@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1838.asp
    profession: Technicien agricole
    site_web: http://www.jeanlassalle.fr
    debut_mandat: 20/06/2007
    nom: Jean Lassalle
    type: depute
  depute_1844:
    fonctions:
      - commission des finances / secrétaire / 
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
    sexe: H
    id_an: 1844
    extras:
      - conférence de la ruralité / membre titulaire
      - comité d'enquête sur le coût et le rendement des services publics / membre titulaire
    adresses:
      - Permanence 5 Rue Roquefort BP 99 46103 Figeac Cedex Téléphone : 05 65 34 12 46 Télécopie : 05 65 34 76 07 
      - Mairie 46130 Bretenoux Téléphone : 05 65 33 81 42 Télécopie : 05 65 39 75 89 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Lot (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Launay
    place_hemicycle: 469
    autresmandats:
      - Maire de Bretenoux, Lot (1231 habitants)
      - Vice-président de la Communauté de communes Cère et Dordogne
    mails:
      - launay.depute@wanadoo.fr
      - jlaunay@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1844.asp
    profession: Inspecteur du Trésor
    site_web: http://www.jeanlaunay.com
    debut_mandat: 20/06/2007
    nom: Jean Launay
    type: depute
  depute_1857:
    place_hemicycle: 334
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Maire de Phalempin, Nord (4615 habitants)
    sexe: H
    id_an: 1857
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1857.asp
    mails:
      - Thierry.LAZARO@wanadoo.fr
      - tlazaro@assemblee-nationale.fr
    adresses:
      - 95 Rue du Général de Gaulle 59133 Phalempin 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chargé de communication
    debut_mandat: 20/06/2007
    nom_de_famille: Lazaro
    nom: Thierry Lazaro
    type: depute
  depute_1866:
    place_hemicycle: 607
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 1866
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1866.asp
    mails:
      - glebris@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 1 Rue du Pladen 29900 Concarneau cedex 
    circonscription: Finistère (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.gilbertlebris.net 
    profession: Commerçant
    debut_mandat: 20/06/2007
    nom_de_famille: Bris
    nom: Gilbert Le Bris
    type: depute
  depute_1871:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1871
    extras:
      - haut comité pour la transparence et l'information sur la sécurité nucléaire / membre titulaire
    adresses:
      - Permanence parlementaire 14 Rue Victor Hugo BP 177 54706 Pont-à-Mousson cedex Téléphone : 03 83 82 13 81 Télécopie : 03 83 82 40 95 
      - Permanence 3 Rue Joffre 54150 Briey Téléphone : 03 82 46 67 33 Télécopie : 03 82 20 97 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meurthe-et-Moselle (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Déaut
    place_hemicycle: 447
    autresmandats:
      - Premier Vice-président du conseil régional (Lorraine)
    mails:
      - jyledeaut@assemblee-nationale.fr
      - jean-yves.le-deaut@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1871.asp
    profession: Professeur d'Université
    site_web: http://www.jyledeaut.fr
    debut_mandat: 20/06/2007
    nom: Jean-Yves Le Déaut
    type: depute
  depute_1874:
    fonctions:
      - assemblée nationale / vice-président / 27/06/2007
      - commission des finances / membre / 
      - délégation chargée des représentants d'intérêts / président / 
      - délégation spéciale chargée de la question des groupes d'intérêt / président / 
      - délégation chargée de l'informatique et des nouvelles technologies / membre / 
      - délégation chargée des groupes d'études et des offices parlementaires / président / 
    sexe: H
    id_an: 1874
    adresses:
      - Permanence 6 Avenue des Combattants 22600 Loudéac Téléphone : 02 96 66 42 63 Télécopie : 02 96 66 42 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côtes-d'Armor (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Fur
    place_hemicycle: 54
    autresmandats:
      - Membre du conseil général (Côtes-d'Armor)
    mails:
      - mlefur@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1874.asp
    profession: Sous-préfet
    site_web: http://www.marclefur.com
    debut_mandat: 20/06/2007
    nom: Marc Le Fur
    type: depute
  depute_1880:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 1880
    extras:
      - haut conseil pour l'avenir de l'assurance maladie / membre titulaire
    adresses:
      - Parti Socialiste 147 Avenue de Choisy 75013 Paris Téléphone : 01 45 86 60 49 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (9ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Guen
    place_hemicycle: 433
    autresmandats:
      - Adjoint au Maire de Paris, Paris (2121291 habitants)
      - Conseiller de Paris
    mails:
      - jmleguen@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1880.asp
    profession: Médecin 
    debut_mandat: 20/06/2007
    nom: Jean-Marie Le Guen
    type: depute
  depute_1883:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 1883
    adresses:
      - Permanence 7 Rue de la Libération 56240 Plouay Téléphone : 02 97 33 19 80 Télécopie : 02 97 33 19 79 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Morbihan (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Nay
    place_hemicycle: 335
    autresmandats:
      - Maire de Plouay, Morbihan (4759 habitants)
    mails:
      - jlenay@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1883.asp
    profession: Horticulteur
    site_web: http://www.jacques-lenay.org
    debut_mandat: 20/06/2007
    nom: Jacques Le Nay
    type: depute
  depute_1886:
    place_hemicycle: 421
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 1886
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1886.asp
    mails:
      - bleroux@assemblee-nationale.fr
      - brunolerouxdepute@yahoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.brunoleroux-blog.org
    profession: Consultant en gestion et management
    debut_mandat: 20/06/2007
    nom_de_famille: Roux
    nom: Bruno Le Roux
    type: depute
  depute_1893:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
      - délégation chargée de la communication et de la presse / questeure, membre / 
      - délégation chargée de l'informatique et des nouvelles technologies / questeure, membre / 
      - délégation chargée de la communication audiovisuelle et de la presse / questeure, membre / 
      - assemblée nationale / questeure / 27/06/2007
    sexe: F
    id_an: 1893
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
      - conseil national du littoral / membre titulaire
    adresses:
      - 6  Place Emile Souvestre 29600 Morlaix Téléphone : 02 98 88 10 09 Télécopie : 02 98 63 44 85 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Finistère (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lebranchu
    place_hemicycle: 500
    autresmandats:
      - Premier Vice-président du conseil régional (Bretagne)
    mails:
      - mlebranchu@assemblee-nationale.fr
      - permanence.lebranchu@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1893.asp
    profession: Vacataire professionnelle à l'Université
    site_web: http://www.lebranchu.fr
    debut_mandat: 20/06/2007
    nom: Marylise Lebranchu
    type: depute
  depute_1911:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1911
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie d'Arques-Cabinet parlementaire Place Roger Salengro BP 60067 Arques 62507 Saint-Omer Cedex Téléphone : 03 21 12 62 30 Télécopie : 03 21 98 80 25 
    circonscription: Pas-de-Calais (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lefait
    place_hemicycle: 513
    autresmandats:
      - Vice-président du conseil général (Pas-de-Calais)
    mails:
      - lefait.michel@wanadoo.fr
      - mlefait@assemblee-nationale.fr
      - ass.nat.lefait.michel@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1911.asp
    profession: Professeur de collège
    site_web: http://michellefait.com  
    debut_mandat: 20/06/2007
    nom: Michel Lefait
    type: depute
  depute_1931:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Conseiller de Paris
    sexe: H
    id_an: 1931
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1931.asp
    mails:
      - plellouche@assemblee-nationale.fr
      - pierre.lellouche@wanadoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire (8e et 9e) 9 Bis Rue de Maubeuge 75009 Paris Téléphone : 01 48 78 24 10 Télécopie : 01 48 78 24 03 
    circonscription: Paris (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Avocat et universitaire
    debut_mandat: 20/06/2007
    nom_de_famille: Lellouche
    nom: Pierre Lellouche
    type: depute
  depute_1936:
    place_hemicycle: 540
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Membre du conseil général (Haute-Garonne)
      - Membre du Conseil municipal de Montesquieu-Volvestre, Haute-Garonne (2314 habitants)
    sexe: H
    id_an: 1936
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1936.asp
    mails:
      - Patrick.LEMASLE@wanadoo.fr
      - plemasle@assemblee-nationale.fr
    adresses:
      - 21 Rue du Faubourg Saint-Germain 31310 Montesquieu-Volvestre Téléphone : 05 61 98 41 93 Télécopie : 05 61 90 52 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Exploitant agricole
    debut_mandat: 20/06/2007
    nom_de_famille: Lemasle
    nom: Patrick Lemasle
    type: depute
  depute_1942:
    fonctions:
      - mission d'information commune sur les prix des carburants dans les dom / membre / 
      - commission des affaires économiques / secrétaire / 
    sexe: H
    id_an: 1942
    extras:
      - conseil supérieur de l'énergie / membre titulaire
    adresses:
      - Hôtel de Ville Place du Général de Gaulle BP 85 61400 Mortagne-au-Perche Téléphone : 02 33 85 11 27 Télécopie : 02 33 25 34 62 
      - Permanence parlementaire 40 Rue Saint-Jean 61300 L'Aigle Téléphone : 02 33 34 79 39 Télécopie : 02 33 25 34 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Orne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lenoir
    place_hemicycle: 257
    autresmandats:
      - Maire de Mortagne-au-Perche, Orne (4506 habitants)
      - Président Communauté de communes du bassin de Mortagne au Perche
    mails:
      - jclenoir@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1942.asp
    profession: Cadre EDF
    debut_mandat: 20/06/2007
    nom: Jean-Claude Lenoir
    type: depute
  depute_1944:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1944
    extras:
      - commission chargée d'examiner les demandes d'autorisation ou de renouvellement d'autorisation des jeux / membre titulaire
    adresses:
      - Mairie Boulevard de la Libération 17340 Châtelaillon-Plage Téléphone : 05 46 30 18 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Charente-Maritime (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Léonard
    place_hemicycle: 206
    autresmandats:
      - Vice-président de la communauté d'agglomération de La Rochelle
      - Maire de Châtelaillon-Plage, Charente-Maritime (5613 habitants)
    mails:
      - jl.leonard@chatelaillonplage.fr
      - jlleonard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1944.asp
    profession: Ingénieur
    site_web: http://www.jeanlouisleonard.com
    debut_mandat: 20/06/2007
    nom: Jean-Louis Léonard
    type: depute
  depute_1946:
    place_hemicycle: 181
    fonctions:
      - mission d'évaluation de la loi n°2005-370 du 22 avril 2005 relative aux droits des malades et à la fin de vie / rapporteur / 
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire d'Antibes, Alpes-Maritimes (72376 habitants)
    sexe: H
    id_an: 1946
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1946.asp
    mails:
      - jaleonetti@assemblee-nationale.fr
    adresses:
      - Mairie Cours Masséna 06600 Antibes Téléphone : 04 92 90 50 05 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-Maritimes (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Praticien hospitalier
    debut_mandat: 20/06/2007
    nom_de_famille: Leonetti
    nom: Jean Leonetti
    type: depute
  depute_1954:
    place_hemicycle: 269
    fonctions:
      - commission des affaires européennes / président / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Vice-président du conseil général (Yvelines)
    sexe: H
    id_an: 1954
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1954.asp
    mails:
      - plequiller@assemblee-nationale.fr
    adresses:
      - Conseil général des Yvelines 2 Place André Mignot 78012 Versailles cedex Téléphone : 01 39 07 76 53 Télécopie : 01 39 07 88 89 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 43 34 Télécopie : 01 40 63 43 43 
    circonscription: Yvelines (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre de banque
    debut_mandat: 20/06/2007
    nom_de_famille: Lequiller
    nom: Pierre Lequiller
    type: depute
  depute_1960:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 1960
    extras:
      - conseil national de l'aménagement et du développement du territoire / membre titulaire
    adresses:
      - Permanence 32    Mail Leclerc 41100 Vendôme Téléphone : 02 54 89 01 72 Télécopie : 02 54 89 01 75 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loir-et-Cher (3ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Leroy
    place_hemicycle: 376
    autresmandats:
      - Président du conseil général (Loir-et-Cher)
    mails:
      - mleroy@assemblee-nationale.fr
      - mleroy.depute@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1960.asp
    profession: Économiste
    debut_mandat: 20/06/2007
    nom: Maurice Leroy
    type: depute
  depute_1977:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 1977
    adresses:
      - 4 Rue Jacques Tourneur BP 90069 57703 Hayange cedex Téléphone : 03 82 84 06 06 Télécopie : 03 82 84 66 88 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Moselle (10ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Liebgott
    place_hemicycle: 551
    autresmandats:
      - Maire de Fameck, Moselle (12635 habitants)
      - Vice-président de la Communauté d'agglomération du Val de Fensch
    mails:
      - mliebgott@assemblee-nationale.fr
      - michel.liebgott@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1977.asp
    profession: Inspecteur des affaires sanitaires et sociales
    site_web: http://www.michel-liebgott.com
    debut_mandat: 20/06/2007
    nom: Michel Liebgott
    type: depute
  depute_1979:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: F
    id_an: 1979
    extras:
      - conseil supérieur du service public ferroviaire / membre titulaire
    adresses:
      - Permanence parlementaire 56 Rue Émile Guichenné BP 621 64006 Pau cedex Téléphone : 05 59 82 20 80 Télécopie : 05 59 82 20 84 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Atlantiques (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lignières-Cassou
    place_hemicycle: 410
    autresmandats:
      - Présidente Communauté d'Agglomération de Pau Pyrénées
      - Maire de Pau, Pyrénées-Atlantiques (81000 habitants)
    mails:
      - martine.lignieres-cassou@wanadoo.fr
      - mlignieres@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1979.asp
    profession: Chargée d'études à la DDE des Pyrénées-Atlantiques
    site_web: http://www.martine-lignieres-cassou.fr/
    debut_mandat: 20/06/2007
    nom: Martine Lignières-Cassou
    type: depute
  depute_1991:
    place_hemicycle: 526
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 1991
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1991.asp
    mails:
      - francois.loncle@wanadoo.fr
      - floncle@assemblee-nationale.fr
    adresses:
      - 17 Rue du Rempart 27400 Louviers Téléphone : 02 32 40 58 80 Télécopie : 02 32 40 45 13 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Eure (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Journaliste
    debut_mandat: 20/06/2007
    nom_de_famille: Loncle
    nom: François Loncle
    type: depute
  depute_1994:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 1994
    extras:
      - conseil de surveillance de l'agence de l'innovation industrielle / membre titulaire
      - observatoire national du service public de l'électricité et du gaz / membre titulaire
      - conseil de surveillance de l'agence française de développement / membre titulaire
    adresses:
      - 5A Rue du Maréchal Foch 67500 Haguenau Téléphone : 03 88 93 63 40 Télécopie : 03 88 93 24 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Loos
    place_hemicycle: 162
    autresmandats:
      - Membre du conseil régional (Alsace)
    mails:
      - francois.loos@yahoo.fr
      - floos@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/1994.asp
    profession: Ingénieur en chef des mines
    debut_mandat: 20/06/2007
    nom: François Loos
    type: depute
  depute_2011:
    fonctions:
      - commission des affaires européennes / membre / 
      - assemblée nationale / secrétaire / 27/06/2007
      - délégation chargée des représentants d'intérêts / membre / 
      - commission des affaires étrangères / membre / 
      - délégation spéciale chargée de la question des groupes d'intérêt / membre / 
      - délégation chargée des groupes d'études et des offices parlementaires / membre / 
    sexe: H
    id_an: 2011
    extras:
      - observatoire national de la sécurité des établissements scolaires et d'enseignement supérieur / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 14 Rue Jean-Raymond Giacosa 06800 Cagnes-sur-Mer Téléphone : 04 93 22 94 44 Télécopie : 04 93 22 96 66 
    circonscription: Alpes-Maritimes (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Luca
    place_hemicycle: 276
    autresmandats:
      - Membre du conseil général (Alpes-Maritimes)
    mails:
      - ll@lionnel-luca.org
      - lluca@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2011.asp
    profession: Professeur d'histoire-géographie
    site_web: http://www.lionnel-luca.org
    debut_mandat: 20/06/2007
    nom: Lionnel Luca
    type: depute
  depute_2045:
    fonctions:
      - commission des lois / secrétaire / 
    sexe: H
    id_an: 2045
    extras:
      - commission nationale consultative des gens du voyage / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville, Cabinet du Maire Rue Calixte Camelle BP 153 33321 Bègles Téléphone : 05 56 49 88 14 Télécopie : 05 56 49 23 79 
    circonscription: Gironde (3ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Mamère
    place_hemicycle: 596
    autresmandats:
      - Maire de Bègles, Gironde (22475 habitants)
    mails:
      - nmamere@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2045.asp
    profession: Journaliste
    site_web: http://www.noelmamere.fr
    debut_mandat: 20/06/2007
    nom: Noël Mamère
    type: depute
  depute_2048:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2048
    extras:
      - conseil d'administration du centre national d'art et de culture georges pompidou / membre titulaire
    adresses:
      - Conseil général de l'Oise 1 Rue Cambry 60000 Beauvais Téléphone : 03 44 06 60 67 Télécopie : 03 44 06 63 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mancel
    place_hemicycle: 280
    autresmandats:
      - Président de la communauté de communes du Pays-de-Thelle
      - Membre du Conseil municipal de Novillers, Oise (315 habitants)
      - Membre du conseil général (Oise)
    mails:
      - jfmancel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2048.asp
    profession: Administrateur civil
    site_web: http://www.jfmancel.com
    debut_mandat: 20/06/2007
    nom: Jean-François Mancel
    type: depute
  depute_2073:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des affaires européennes / vice-président / 
      - commission des lois / membre / 
    sexe: H
    id_an: 2073
    extras:
      - conseil national de sécurité civile / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 91 25 Télécopie : 01 40 63 91 37 
      - 82 Avenue Charles de Gaulle 84100 Orange Téléphone : 04 90 11 00 00 Télécopie : 04 90 11 06 81 
    circonscription: Vaucluse (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mariani
    place_hemicycle: 93
    autresmandats:
      - Membre du conseil régional (Provence-Alpes-Côte-d'Azur)
    mails:
      - tmariani@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2073.asp
    profession: Cadre
    site_web: http://www.thierrymariani.fr
    debut_mandat: 20/06/2007
    nom: Thierry Mariani
    type: depute
  depute_2075:
    place_hemicycle: 591
    fonctions:
      - mission d'information commune sur les prix des carburants dans les dom / membre / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Président du conseil régional (Martinique)
    sexe: H
    id_an: 2075
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2075.asp
    mails:
      - amarie@assemblee-nationale.fr
    adresses:
      - Mairie 97211 Rivière-Pilote Téléphone : 05 96 62 60 03 Télécopie : 05 96 62 73 65 
      - Circonscription 12, Rue Paul Langevin 97228 Saint-Luce Téléphone : 05 96 62 30 62 Télécopie : 05 96 62 29 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Martinique (4ème)
    groupe:
      - gauche démocrate et républicaine / membre
    profession: Professeur de mathématiques
    debut_mandat: 20/06/2007
    nom_de_famille: Marie-Jeanne
    nom: Alfred Marie-Jeanne
    type: depute
  depute_2083:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / rapporteur / 
      - commission des finances / membre / 
    sexe: H
    id_an: 2083
    extras:
      - comité d'orientation du centre d'analyse stratégique / membre titulaire
      - conseil supérieur de la coopération / membre titulaire
      - conseil d'administration du fonds pour le développement de l'intermodalité dans les transports / membre titulaire
      - conseil national de l'information statistique / membre titulaire
    adresses:
      - Permanence 5 Rue Paul Pons 26400 Crest Téléphone : 04 75 76 71 34 Télécopie : 04 75 25 44 56 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Drôme (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mariton
    place_hemicycle: 78
    autresmandats:
      - Maire de Crest, Drôme (7744 habitants)
    mails:
      - hmariton@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2083.asp
    profession: Ingénieur en chef des mines
    site_web: http://www.herve-mariton.net
    debut_mandat: 20/06/2007
    nom: Hervé Mariton
    type: depute
  depute_2086:
    place_hemicycle: 18
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Maire d'Étampes, Essonne (21839 habitants)
    sexe: H
    id_an: 2086
    mails:
      - depute@franckmarlin.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2086.asp
    circonscription: Essonne (2ème)
    adresses:
      - Hôtel de Ville BP 109 91152 Étampes cedex Téléphone : 01 69 92 68 91 Télécopie : 01 69 92 68 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    groupe:
      - union pour un mouvement populaire / apparenté
    debut_mandat: 20/06/2007
    nom_de_famille: Marlin
    nom: Franck Marlin
    type: depute
  depute_2098:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2098
    extras:
      - conseil de modération et de prévention / membre titulaire
    adresses:
      - 15 Rue Jean Moët 51200 Épernay Téléphone : 03 26 59 30 04 Télécopie : 03 26 59 99 81 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Marne (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Martin
    place_hemicycle: 11
    autresmandats:
      - Adjoint au Maire de Cumières, Marne (861 habitants)
      - Vice-président de la communauté de communes d'Epernay Pays de Champagne
    mails:
      - pamartin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2098.asp
    profession: Viticulteur
    debut_mandat: 20/06/2007
    nom: Philippe Armand Martin
    type: depute
  depute_2099:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2099
    extras:
      - conseil consultatif de l'internet / membre titulaire
      - commission nationale consultative des gens du voyage / membre titulaire
      - conseil supérieur de l'énergie / membre suppléant
    adresses:
      - Cabinet parlementaire 4 Place de la Paix BP 119 41203 Romorantin-Lanthenay cedex Téléphone : 02 54 76 76 53 Télécopie : 02 54 76 44 66 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loir-et-Cher (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Martin-Lalande
    place_hemicycle: 125
    autresmandats:
      - Membre du conseil général (Loir-et-Cher)
    mails:
      - pmartin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2099.asp
    profession: Cadre administratif
    debut_mandat: 20/06/2007
    nom: Patrice Martin-Lalande
    type: depute
  depute_2102:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: F
    id_an: 2102
    extras:
      - commission de surveillance et de contrôle des publications destinées à l'enfance et à l'adolescence / membre suppléante
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 72 76 Télécopie : 01 40 63 78 24 
      - Secrétariat parlementaire 24 Rue Carnot 05000 Gap Téléphone : 04 92 52 38 72 Télécopie : 04 92 56 23 84 
    circonscription: Hautes-Alpes (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Martinez
    place_hemicycle: 199
    autresmandats:
      - Membre du Conseil municipal de Laragne-Montéglin, Hautes-Alpes (3296 habitants)
    mails:
      - henriette.martinez@wanadoo.fr
      - hmartinez@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2102.asp
    profession: Professeur certifié
    site_web: http://www.henriettemartinez.com
    debut_mandat: 20/06/2007
    nom: Henriette Martinez
    type: depute
  depute_210741:
    place_hemicycle: 527
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Vice-président du conseil général (Pas-de-Calais)
    sexe: H
    id_an: 210741
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/210741.asp
    mails:
      - Jean-Claude.Leroy9@wanadoo.fr
      - jcleroy@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 2 Place Jean Jaurès BP 45 62380 Lumbres Téléphone : 03 21 38 76 76 Télécopie : 03 21 38 76 78 
    circonscription: Pas-de-Calais (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Attaché territorial
    debut_mandat: 20/06/2007
    nom_de_famille: Leroy
    nom: Jean-Claude Leroy
    type: depute
  depute_2107:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 2107
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence  16 Avenue du Cep 78300 Poissy Téléphone : 01 30 74 43 69 Télécopie : 01 39 79 42 24 
    circonscription: Yvelines (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Masdeu-Arus
    place_hemicycle: 266
    autresmandats:
      - Membre du Conseil municipal de Poissy, Yvelines (35841 habitants)
    mails:
      - jmasdeu@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2107.asp
    profession: Ingénieur conseil
    site_web: http://www.jmasdeu-arus.com
    debut_mandat: 20/06/2007
    nom: Jacques Masdeu-Arus
    type: depute
  depute_211169:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 211169
    adresses:
      - Mairie 177 Avenue Gabriel Péri 92230 Gennevilliers Téléphone : 01 40 85 62 30 Télécopie : 01 47 99 07 56 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 88 
    circonscription: Hauts-de-Seine (1ère)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Muzeau
    place_hemicycle: 584
    autresmandats:
      - Premier adjoint de Gennevilliers, Hauts-de-Seine (42612 habitants)
    mails:
      - rmuzeau@assemblee-nationale.fr
      - r.muzeau@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/211169.asp
    profession: Ajusteur-outilleur
    site_web: http://www.roland-muzeau.org
    debut_mandat: 20/06/2007
    nom: Roland Muzeau
    type: depute
  depute_2124:
    fonctions:
      - commission des finances / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
    sexe: H
    id_an: 2124
    extras:
      - conseil supérieur des prestations sociales agricoles / membre titulaire
      - comité de surveillance du fonds de solidarité vieillesse / membre titulaire
    adresses:
      - Mairie Château Saint-Louis 10340 Les Riceys Téléphone : 03 25 29 30 32 Télécopie : 03 25 29 72 09 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 2 Rue des Anciennes Tanneries 10000 Troyes Téléphone : 03 25 41 86 87 Télécopie : 03 25 41 86 88 
    circonscription: Aube (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mathis
    place_hemicycle: 220
    autresmandats:
      - Vice-président du conseil général (Aube)
      - Maire des Riceys, Aube (1376 habitants)
    mails:
      - jcmathis@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2124.asp
    profession: Directeur de société
    debut_mandat: 20/06/2007
    nom: Jean-Claude Mathis
    type: depute
  depute_2126:
    fonctions:
      - commission des affaires étrangères / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / vice-président / 
    sexe: H
    id_an: 2126
    extras:
      - conseil d'administration de l'institut national de l'audiovisuel (ina) / membre titulaire
    adresses:
      - Hôtel de Ville 18  Rue Carnot BP 188 71307 Montceau-les-Mines cedex Téléphone : 03 85 67 68 30 Télécopie : 03 85 67 68 32 
      - Permanence parlementaire 4 Rue Carnot BP 202 71308 Montceau-les-Mines cedex Téléphone : 03 85 57 03 88 Télécopie : 03 85 58 69 47 
      - Communauté urbaine Le Creusot Monceau Château de la Verrerie BP 69 71206 Le Creusot cedex Télécopie : 03 85 56 38 51 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Mathus
    place_hemicycle: 524
    autresmandats:
      - Maire de Montceau-les-Mines, Saône-et-Loire (20632 habitants)
    mails:
      - mathus.didier@wanadoo.fr
      - dmathus@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2126.asp
    profession: Enseignant
    site_web: http://www.didiermathus.com
    debut_mandat: 20/06/2007
    nom: Didier Mathus
    type: depute
  depute_2148:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des affaires sociales / président / 
    sexe: H
    id_an: 2148
    extras:
      - conseil d'orientation des finances publiques / membre titulaire
      - haut conseil pour l'avenir de l'assurance maladie / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie BP 70627 35506 Vitré cedex Téléphone : 02 99 75 07 28 
    circonscription: Ille-et-Vilaine (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Méhaignerie
    place_hemicycle: 186
    autresmandats:
      - Président de la communauté d'agglomération de Vitré communauté
      - Maire de Vitré, Ille-et-Vilaine (15282 habitants)
    mails:
      - pmehaignerie@assemblee-nationale.fr
      - pmehaign@club-internet.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2148.asp
    profession: Ingénieur du génie rural et des eaux et forêts
    site_web: http://www.pierre-mehaignerie.org
    debut_mandat: 20/06/2007
    nom: Pierre Méhaignerie
    type: depute
  depute_216574:
    place_hemicycle: 399
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Pfastatt, Haut-Rhin (8500 habitants)
    sexe: H
    id_an: 216574
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/216574.asp
    mails:
      - fhillmeyer@assemblee-nationale.fr
      - FRANCIS.HILLMEYER@wanadoo.fr
    adresses:
      - 128 Rue de la République 68120 Pfastatt Téléphone : 03 89 53 59 92 Télécopie : 03 89 53 57 38 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (6ème)
    groupe:
      - nouveau centre / membre
    profession: Journaliste reporter-photographe
    debut_mandat: 20/06/2007
    nom_de_famille: Hillmeyer
    nom: Francis Hillmeyer
    type: depute
  depute_2181:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 2181
    extras:
      - haut conseil du secteur public / membre titulaire
    adresses:
      - Permanence 36 Avenue Archon-Despérouses 63200 Riom Téléphone : 04 73 38 66 03 Télécopie : 04 73 38 66 45 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Puy-de-Dôme (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Michel
    place_hemicycle: 445
    autresmandats:
      - Maire de Lapeyrouse, Puy-de-Dôme (587 habitants)
    mails:
      - jean.michel10@wanadoo.fr
      - jmichel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2181.asp
    profession: Avocat
    debut_mandat: 20/06/2007
    nom: Jean Michel
    type: depute
  depute_2189:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission des finances) de la mission d'évaluation et de contrôle (commission des finances) / (président / 
      - commission des finances / président / 
    sexe: H
    id_an: 2189
    extras:
      - conseil d'orientation des finances publiques / membre titulaire
    adresses:
      - 20 Avenue de la Houille Blanche 38170 Seyssinet-Pariset Téléphone : 04 76 70 15 15 Télécopie : 04 76 70 15 16 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Migaud
    place_hemicycle: 514
    autresmandats:
      - Maire de Seyssins, Isère (6850 habitants)
      - Président de la communauté d'agglomération Grenoble-Alpes Métropole
    mails:
      - dmigaud@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2189.asp
    profession: Juriste
    site_web: http://www.didiermigaud.fr
    debut_mandat: 20/06/2007
    nom: Didier Migaud
    type: depute
  depute_2191:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2191
    adresses:
      - BP 11 77630 Barbizon Téléphone : 01 60 66 42 58 Télécopie : 01 60 66 42 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Autre téléphone : 01 40 63 67 97 Autre télécopie : 01 40 63 99 79  Jean-claude.MIGNON@wanadoo.fr
    circonscription: Seine-et-Marne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mignon
    place_hemicycle: 27
    autresmandats:
      - Maire de Dammarie-les-Lys, Seine-et-Marne (20659 habitants)
    mails:
      - jcmignon@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2191.asp
    profession: Ancien chef d'entreprise
    site_web: http://www.jean-claude-mignon.net
    debut_mandat: 20/06/2007
    nom: Jean-Claude Mignon
    type: depute
  depute_2224:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 2224
    adresses:
      - 9 Rue des Dôdanes 71500 Louhans Téléphone : 03 85 75 76 77 Télécopie : 03 85 75 76 70 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Montebourg
    place_hemicycle: 503
    autresmandats:
      - Président du conseil général (Saône-et-Loire)
    mails:
      - amontebourg@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2224.asp
    profession: Avocat 
    site_web: http://www.arnaudmontebourg.fr
    debut_mandat: 20/06/2007
    nom: Arnaud Montebourg
    type: depute
  depute_2229:
    fonctions:
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / coprésident / 
      - commission des affaires sociales / vice-président / 
      - mission d'information commune sur les exonérations sociales / membre / 
    sexe: H
    id_an: 2229
    extras:
      - conseil de surveillance de la caisse nationale de l'assurance maladie des travailleurs salariés / membre titulaire
      - conseil d'administration de la société nationale de programme "france 2" / membre titulaire
      - conseil de modération et de prévention / membre titulaire
      - conseil de surveillance de l'agence centrale des organismes de sécurité sociale / membre titulaire
      - commission des comptes de la sécurité sociale / membre titulaire
      - comité national de l'organisation sanitaire et sociale / membre titulaire
    adresses:
      - Permanence parlementaire 2  Rue de la Procession 78100 Saint-Germain-en-Laye Téléphone : 01 34 51 20 20 Télécopie : 01 39 73 68 74 
      - Mairie Place Charles de Gaulle 78240 Chambourcy Téléphone : 01 39 22 31 31 Télécopie : 01 39 22 31 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yvelines (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Morange
    place_hemicycle: 332
    autresmandats:
      - Maire de Chambourcy, Yvelines (5077 habitants)
    mails:
      - pmorange@assemblee-nationale.fr
      - pierre.morange@noos.fr
      - cabinet@chambourcy.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2229.asp
    profession: Médecin généraliste
    site_web: http://www.pierre-morange.fr
    debut_mandat: 20/06/2007
    nom: Pierre Morange
    type: depute
  depute_2237:
    place_hemicycle: 243
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Membre du conseil général (Deux-Sèvres)
    sexe: H
    id_an: 2237
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2237.asp
    mails:
      - jm.morisset@cg79.fr
      - jmmorisset@assemblee-nationale.fr
    adresses:
      - La Cointrie 79310 Saint-Pardoux Téléphone : 05 49 64 23 22 Télécopie : 05 49 63 32 38 
      - Conseil général Place Denfert-Rochereau BP 351 79021 Niort cedex Téléphone : 05 49 06 79 82 Télécopie : 05 49 06 77 32 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Deux-Sèvres (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur informatique
    debut_mandat: 20/06/2007
    nom_de_famille: Morisset
    nom: Jean-Marie Morisset
    type: depute
  depute_223837:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 223837
    extras:
      - conseil d'administration de la société nationale de programme radio-france / membre titulaire
    adresses:
      - Mairie, Cabinet du Maire Place Bernard Cornut-Gentille BP 140 06406 Cannes cedex 
      - Maison du Mouvement 19  Place du Marché Forville 06400 Cannes Téléphone : 04 93 68 08 12 Télécopie : 04 93 68 39 10 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-Maritimes (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Brochand
    place_hemicycle: 103
    autresmandats:
      - Maire de Cannes, Alpes-Maritimes (67304 habitants)
    mails:
      - bbrochand@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/223837.asp
    profession: Cadre du secteur privé retraité
    site_web: http://www.bernard-brochand.com
    debut_mandat: 20/06/2007
    nom: Bernard Brochand
    type: depute
  depute_2240:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2240
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 51 Avenue des Allies 25200 Montbéliard Téléphone : 03 81 32 31 69 Télécopie : 03 81 32 31 67 
    circonscription: Doubs (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Moscovici
    place_hemicycle: 430
    autresmandats:
      - Membre du Conseil municipal de Valentigney, Doubs (12484 habitants)
      - Président de la communauté d'agglomération du Pays-de-Montbéliard
    mails:
      - pmoscovici@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2240.asp
    profession: Conseiller maître à la cour des comptes
    site_web: http://moscovici.typepad.fr/blognational
    debut_mandat: 20/06/2007
    nom: Pierre Moscovici
    type: depute
  depute_2242:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 2242
    extras:
      - conseil d'orientation de l'observatoire national des zones urbaines sensibles / membre titulaire
    adresses:
      - Permanence 23 Rue Denis Roy 95100 Argenteuil Téléphone : 01 39 61 50 81 Télécopie : 01 39 47 99 37 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mothron
    place_hemicycle: 89
    autresmandats:
      - Membre du Conseil municipal d'Argenteuil, Val-d'Oise (94019 habitants)
    mails:
      - gmothron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2242.asp
    profession: Chef des ventes
    site_web: http://www.georges-mothron.fr
    debut_mandat: 20/06/2007
    nom: Georges Mothron
    type: depute
  depute_2250:
    place_hemicycle: 43
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Membre du conseil général (Isère)
      - Maire de Crémieu, Isère (3169 habitants)
    sexe: H
    id_an: 2250
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2250.asp
    mails:
      - moyne-bressand.alain@wanadoo.fr
      - amoyne@assemblee-nationale.fr
    adresses:
      - Mairie 38460 Crémieu Téléphone : 04 74 90 70 92 Télécopie : 04 74 90 88 86 
      - Secrétariat parlementaire Place du 8 mai 1945 38460 Crémieu Téléphone : 04 74 90 74 18 Télécopie : 04 74 90 83 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chef d'entreprise
    debut_mandat: 20/06/2007
    nom_de_famille: Moyne-Bressand
    nom: Alain Moyne-Bressand
    type: depute
  depute_2256:
    fonctions:
      - commission des affaires étrangères / vice-président / 
    sexe: H
    id_an: 2256
    extras:
      - conseil de surveillance de l'agence française de développement / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Fédération UMP 39 Rue Sainte-Cécile 13005 Marseille Téléphone : 04 91 25 62 61 Télécopie : 04 91 80 46 46 
    circonscription: Bouches-du-Rhône (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Muselier
    place_hemicycle: 96
    autresmandats:
      - Premier vice-président de la communauté urbaine Marseille Provence Métropole
      - Membre du Conseil municipal de Marseille 3ème secteur, Bouches-du-Rhône (798021 habitants)
    mails:
      - rmuselier@assemblee-nationale.fr
      - muselier.ump@online.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2256.asp
    profession: Médecin coordonnateur d'un établissement hospitalier privé
    site_web: http://www.renaud-muselier.com
    debut_mandat: 20/06/2007
    nom: Renaud Muselier
    type: depute
  depute_2257:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2257
    adresses:
      - Permanence 36 Avenue de la République 78500 Sartrouville Téléphone : 01 39 13 93 93 
      - Mairie 48 Avenue de Longueil 78600 Maisons-Laffitte Téléphone : 01 34 93 12 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yvelines (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Myard
    place_hemicycle: 292
    autresmandats:
      - Maire de Maisons-Laffitte, Yvelines (21856 habitants)
    mails:
      - jmyard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2257.asp
    profession: Conseiller des affaires étrangères
    site_web: http://www.jacques-myard.org
    debut_mandat: 20/06/2007
    nom: Jacques Myard
    type: depute
  depute_2265:
    place_hemicycle: 352
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Brive-la-Gaillarde, Corrèze (49139 habitants)
    sexe: H
    id_an: 2265
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2265.asp
    mails:
      - pnauche@assemblee-nationale.fr
      - permanence.nauche@orange.fr
    adresses:
      - Permanence parlementaire 2 Rue du maréchal Brune 19100 Brive la Gaillarde Téléphone : 05 55 17 02 86 Télécopie : 05 55 17 03 53 
      - Mairie de Brive Place de l'Hôtel de Ville BP 433 19312 Brive cedex Téléphone : 05 55 18 17 63 Télécopie : 05 55 18 15 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Corrèze (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Médecin hospitalier
    debut_mandat: 20/06/2007
    nom_de_famille: Nauche
    nom: Philippe Nauche
    type: depute
  depute_2269:
    fonctions:
      - commission des finances / membre / 
      - délégation chargée de la communication et de la presse / membre / 
      - assemblée nationale / secrétaire / 01/10/2008
      - délégation chargée de l'informatique et des nouvelles technologies / membre / 
    sexe: H
    id_an: 2269
    adresses:
      - 1 Quai du Gravier BP 40 09201 Saint-Girons cedex Téléphone : 05 61 04 64 64 Télécopie : 05 61 04 65 65 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ariège (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Nayrou
    place_hemicycle: 544
    autresmandats:
      - Membre du conseil général (Ariège)
    mails:
      - hnayrou@assemblee-nationale.fr
      - henri.nayrou@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2269.asp
    profession: Journaliste
    site_web: http://www.henrinayrou.com
    debut_mandat: 20/06/2007
    nom: Henri Nayrou
    type: depute
  depute_226:
    fonctions:
      - commission des affaires économiques / membre / 
      - mission d'information commune sur l'évaluation des dispositifs fiscaux d'encouragement à l'investissement locatif / membre / 
    sexe: H
    id_an: 226
    extras:
      - conseil national de l'habitat / membre titulaire
    adresses:
      - Permanence parlementaire 102 Boulevard Blossac 86100 Châtellerault Téléphone : 05 49 02 15 75 Télécopie : 05 49 02 15 76 
      - Cabinet du Maire 78 Boulevard Blossac BP619 86106 Châtellerault cedex 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vienne (4ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Abelin
    place_hemicycle: 385
    autresmandats:
      - Maire de Châtellerault, Vienne (34126 habitants)
      - Président de la communauté d'agglomération du Pays Châtelleraudais
    mails:
      - jpabelin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/226.asp
    profession: Directeur-adjoint de service à la Banque de France
    site_web: http://www.jpabelin.com
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Abelin
    type: depute
  depute_2272:
    place_hemicycle: 522
    fonctions:
      - commission des affaires étrangères / membre / 
      - délégation chargée d'examiner la recevabilité des propositions de loi / président / 
      - assemblée nationale / vice-président / 01/10/2008
      - délégation chargée de l'informatique et des nouvelles technologies / membre / 
    autresmandats:
      - Maire de Beauregard-l'Évêque, Puy-de-Dôme (1158 habitants)
      - Membre du conseil général (Puy-de-Dôme)
    sexe: H
    id_an: 2272
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2272.asp
    mails:
      - aneri@assemblee-nationale.fr
    adresses:
      - 100 Avenue Léon Blum 63000 Clermont-Ferrand Téléphone : 04 73 26 01 85 Télécopie : 04 73 27 78 91 
      - Mairie 63116 Beauregard-l'Évêque Téléphone : 04 73 68 16 03 Télécopie : 04 73 68 07 10 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Puy-de-Dôme (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Retraité de l'Education nationale
    debut_mandat: 20/06/2007
    nom_de_famille: Néri
    nom: Alain Néri
    type: depute
  depute_2273:
    place_hemicycle: 336
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Maire de Paray-le-Monial, Saône-et-Loire (9194 habitants)
    sexe: H
    id_an: 2273
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2273.asp
    mails:
      - jmnesme@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville 13 Place de l'Hôtel de ville 71600 Paray-le-Monial Téléphone : 03 85 81 95 14 Télécopie : 03 85 81 19 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre consulaire
    debut_mandat: 20/06/2007
    nom_de_famille: Nesme
    nom: Jean-Marc Nesme
    type: depute
  depute_2277:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2277
    adresses:
      - 4 Rue Molière BP 273 42301 Roanne cedex Téléphone : 04 77 70 98 98 Télécopie : 04 77 70 93 10 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Nicolin
    place_hemicycle: 265
    autresmandats:
      - Membre du Conseil municipal de Roanne, Loire (38887 habitants)
    mails:
      - ynicolin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2277.asp
    profession: Gestionnaire
    site_web: http://www.yvesnicolin.fr
    debut_mandat: 20/06/2007
    nom: Yves Nicolin
    type: depute
  depute_2295:
    fonctions:
      - mission d'information commune sur les prix des carburants dans les dom / président / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des affaires économiques / président / 
    sexe: H
    id_an: 2295
    adresses:
      - Mairie 92501 Rueil-Malmaison Téléphone : 01 47 32 66 29 Télécopie : 01 47 32 67 84 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hauts-de-Seine (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ollier
    place_hemicycle: 180
    autresmandats:
      - Maire de Rueil-Malmaison, Hauts-de-Seine (73469 habitants)
    mails:
      - pollier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2295.asp
    profession: Cadre de société
    site_web: http://www.patrick-ollier.com
    debut_mandat: 20/06/2007
    nom: Patrick Ollier
    type: depute
  depute_230329:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 230329
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (13ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lamour
    place_hemicycle: 101
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Conseiller de Paris
    mails:
      - jflamour@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/230329.asp
    profession: Kinésithérapeute
    site_web: http://www.jeanfrancoislamour.fr
    debut_mandat: 20/06/2007
    nom: Jean-François Lamour
    type: depute
  depute_230:
    place_hemicycle: 77
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / président / 
      - assemblée nationale / président / 26/06/2007
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Premier vice-président de la communauté d'agglomération d'Annecy
      - Maire d'Annecy-le-Vieux, Haute-Savoie (18885 habitants)
    sexe: H
    id_an: 230
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/230.asp
    mails:
      - baccoyer@assemblee-nationale.fr
      - bernard.accoyer@wanadoo.fr
    adresses:
      - 49 Avenue de Genève 74000 Annecy Téléphone : 04 50 57 57 62 
      - Mairie 74940 Annecy-le-Vieux Téléphone : 04 50 23 86 33 Télécopie : 04 50 27 66 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Savoie (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin ORL
    debut_mandat: 20/06/2007
    nom_de_famille: Accoyer
    nom: Bernard Accoyer
    type: depute
  depute_2317:
    place_hemicycle: 499
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Noisy-le-Grand, Seine-Saint-Denis (58217 habitants)
    sexe: H
    id_an: 2317
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2317.asp
    mails:
      - mpajon@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville Place de la Libération BP 49 93161 Noisy-le-Grand cedex Téléphone : 01 45 92 76 67 Téléphone : 01 45 92 76 90 Télécopie : 01 43 05 27 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 69 86 Télécopie : 01 40 63 91 58 
    circonscription: Seine-Saint-Denis (13ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Maître de conférence en économie (Paris I)
    debut_mandat: 20/06/2007
    nom_de_famille: Pajon
    nom: Michel Pajon
    type: depute
  depute_2319:
    place_hemicycle: 177
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Conseillère de Paris
    sexe: F
    id_an: 2319
    extras:
      - commission nationale pour l'éducation, la science et la culture ( unesco ) / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2319.asp
    mails:
      - fdepanafieu@assemblee-nationale.fr
    adresses:
      - 74 Rue Pierre Demours 75017 Paris Téléphone : 01 43 80 19 10 Télécopie : 01 43 80 24 11 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 66 03 Télécopie : 01 40 63 66 35 
    circonscription: Paris (16ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Panafieu
    nom: Françoise de Panafieu
    type: depute
  depute_2338:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 2338
    extras:
      - commission du dividende numérique / membre titulaire
      - commission nationale des comptes de la formation professionnelle / membre titulaire
      - conseil d'administration de l'ecole nationale d'administration / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 11 
      - Permanence parlementaire 1 Rue des Teuraux 58140 Lormes Téléphone : 03 86 22 89 50 Télécopie : 03 86 22 58 32 
    circonscription: Nièvre (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Paul
    place_hemicycle: 502
    autresmandats:
      - Membre de la Communauté de communes des Portes du Morvan
      - Vice-président du conseil régional (Bourgogne)
      - Membre du Conseil municipal de Lormes, Nièvre (1396 habitants)
    mails:
      - christian.paul@wanadoo.fr
      - cpaul@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2338.asp
    profession: Administrateur civil
    site_web: http://www.christianpaul.fr
    debut_mandat: 20/06/2007
    nom: Christian Paul
    type: depute
  depute_2339:
    fonctions:
      - commission des affaires économiques / secrétaire / 
    sexe: H
    id_an: 2339
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
    adresses:
      - 12 Rue Michel Gautier 76600 Le Havre Téléphone : 02 35 53 05 79 Télécopie : 02 35 53 66 91 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (8ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Paul
    place_hemicycle: 588
    autresmandats:
      - Membre du Conseil municipal du Havre, Seine-Maritime (190590 habitants)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2339.asp
    mails:
      - an.dpaul@wanadoo.fr
    site_web: http://www.danielpaul-lehavre.org
    profession: Instituteur
    debut_mandat: 20/06/2007
    nom: Daniel Paul
    type: depute
  depute_2343:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2343
    extras:
      - comité de surveillance de l'établissement de gestion du fonds de financement des prestations sociales des non-salariés agricoles / membre titulaire
      - comité national de l'eau / membre titulaire
      - conseil supérieur des prestations sociales agricoles / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 14 Place de la Bouquerie BP 75 24202 Sarlat cedex Téléphone : 05 53 31 31 81 Télécopie : 05 53 31 31 84 
    circonscription: Dordogne (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Peiro
    place_hemicycle: 444
    autresmandats:
      - Maire de Castelnaud-la-Chapelle, Dordogne (424 habitants)
      - Membre du conseil général (Dordogne)
    mails:
      - gpeiro@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2343.asp
    profession: Instituteur
    site_web: http://germinal-peiro.com
    debut_mandat: 20/06/2007
    nom: Germinal Peiro
    type: depute
  depute_2345:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2345
    extras:
      - comité des finances locales / membre titulaire
      - conseil d'orientation pour la prévention des risques naturels majeurs / membre titulaire
    adresses:
      - Hôtel de Ville 39000 Lons-le-Saunier Téléphone : 03 84 47 88 31 Télécopie : 03 84 47 88 96 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Jura (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Pélissard
    place_hemicycle: 84
    autresmandats:
      - Président de la communauté de communes du Bassin-de-Lons-le-Saunier
      - Maire de Lons-le-Saunier, Jura (18483 habitants)
    mails:
      - jacques.pelissard@ville-lons-le-saunier.fr
      - jpelissard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2345.asp
    profession: Avocat
    debut_mandat: 20/06/2007
    nom: Jacques Pélissard
    type: depute
  depute_2357:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2357
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 91 22 Télécopie : 01 40 63 91 41 
      - Permanence 116 Rue Cuvier 69006 Lyon  Téléphone : 04 78 24 41 13 Télécopie : 04 78 24 23 30 
    circonscription: Rhône (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Perben
    place_hemicycle: 83
    autresmandats:
      - Vice-président du conseil général (Rhône)
    mails:
      - dperben@assemblee-nationale.fr
      - contact@perben.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2357.asp
    profession: Sous-préfet
    site_web: http://www.perben.com
    debut_mandat: 20/06/2007
    nom: Dominique Perben
    type: depute
  depute_2365:
    place_hemicycle: 516
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Membre du Conseil municipal de Carcassonne, Aude (43950 habitants)
    sexe: H
    id_an: 2365
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2365.asp
    mails:
      - jean-claude.perez@wanadoo.fr
      - jcperez@assemblee-nationale.fr
    adresses:
      - 2 Rue Barbès BP 158 11004 Carcassonne cedex Téléphone : 04 68 47 49 28 Télécopie : 04 68 47 43 88 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 74 53 Télécopie : 01 40 63 79 09 
    circonscription: Aude (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Secrétaire de mairie
    debut_mandat: 20/06/2007
    nom_de_famille: Perez
    nom: Jean-Claude Perez
    type: depute
  depute_236:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 236
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hauts-de-Seine (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Aeschlimann
    place_hemicycle: 204
    autresmandats:
      - Membre du Conseil municipal d'Asnières-sur-Seine, Hauts-de-Seine (75794 habitants)
    mails:
      - maeschlimann@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/236.asp
    profession: Maître de conférences à l'IEP-Paris
    site_web: http://www.manuel-aeschlimann.fr
    debut_mandat: 20/06/2007
    nom: Manuel Aeschlimann
    type: depute
  depute_2371:
    place_hemicycle: 428
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
      - délégation chargée de la communication audiovisuelle et de la presse / membre / 
    autresmandats:
      - Présidente du conseil général (Haute-Vienne)
    sexe: F
    id_an: 2371
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2371.asp
    mails:
      - mfperol@assemblee-nationale.fr
      - mf.peroldumont@wanadoo.fr
    adresses:
      - Conseil général 43 Avenue de la Libération 87000 Limoges Téléphone : 05 55 45 10 49 Télécopie : 05 55 79 57 81 
      - BP 262 87007 Limoges cedex 1 Téléphone : 05 55 10 18 33 Télécopie : 05 55 10 18 42 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Vienne (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur de collège (en détachement depuis 1997)
    debut_mandat: 20/06/2007
    nom_de_famille: Pérol-Dumont
    nom: Marie-Françoise Pérol-Dumont
    type: depute
  depute_2374:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 2374
    extras:
      - comité de l'initiative française pour les récifs coralliens / membre titulaire
    adresses:
      - 43 Rue du 24 Février BP 88 79003 Niort cedex Téléphone : 05 49 77 29 40 Télécopie : 05 49 77 29 44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Deux-Sèvres (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Gaillard
    place_hemicycle: 534
    autresmandats:
      - Maire de Niort, Deux-Sèvres (56663 habitants)
    mails:
      - ggaillard@assemblee-nationale.fr
      - deputee@genevieve-gaillard.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2374.asp
    profession: Vétérinaire
    site_web: http://www.genevieve-gaillard.com
    debut_mandat: 20/06/2007
    nom: Geneviève Gaillard
    type: depute
  depute_2377:
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - assemblée nationale / secrétaire / 27/06/2007
      - commission des affaires sociales / vice-président / 
    sexe: H
    id_an: 2377
    extras:
      - comité national d'évaluation des dispositifs expérimentaux d'aide aux personnes âgées / membre titulaire
      - commission des comptes de la sécurité sociale / membre titulaire
      - conseil national du tourisme / membre titulaire
    adresses:
      - Permanence parlementaire 227 Boulevard Gambetta 69400 Villefranche-sur-Saône Téléphone : 04 74 68 07 44 Télécopie : 04 74 68 21 57 
      - Hôtel de ville Rue de la Paix 69400 Villefranche-sur-Saône Téléphone :  Téléphone : 04 74 62 60 12 Télécopie : 04 74 62 60 92 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Perrut
    place_hemicycle: 203
    autresmandats:
      - Maire de Villefranche-sur-Saône, Rhône (34893 habitants)
      - Vice-président de la communauté d'agglomération de Villefranche-sur-Saône
    mails:
      - bperrut@wanadoo.fr
      - bperrut@villefranche.net
      - bperrut@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2377.asp
    profession: Avocat
    site_web: http://www.bernardperrut.fr
    debut_mandat: 20/06/2007
    nom: Bernard Perrut
    type: depute
  depute_2421:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 2421
    extras:
      - conseil national de l'enseignement supérieur privé / membre titulaire
      - conseil d'administration de l'office français de protection des réfugiés et du du conseil d'administration de l'office français de protection des réfugiés et apatrides  / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yvelines (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Pinte
    place_hemicycle: 329
    mails:
      - epinte@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2421.asp
    profession: Cadre d'un établissement public
    site_web: http://www.etiennepinte.com
    debut_mandat: 20/06/2007
    nom: Étienne Pinte
    type: depute
  depute_2424:
    place_hemicycle: 338
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Membre du conseil général (Val-de-Marne)
      - Maire de Saint-Maur-des-Fossés, Val-de-Marne (72955 habitants)
    sexe: H
    id_an: 2424
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2424.asp
    mails:
      - hplagnol@assemblee-nationale.fr
    adresses:
      - 37 Avenue Joffre 94100 Saint Maur des Fossés 
      - Hôtel de ville Place Charles de Gaulle 94100 Saint Maur des Fossés Téléphone : 01 45 11 65 13 
      - Conseil général du Val de Marne 21 Avenue du Général de Gaulle Hôtel du Département 94011 Créteil cedex Téléphone : 01 43 99 71 47 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Conseiller d'État - Professeur associé à Paris Dauphine
    debut_mandat: 20/06/2007
    nom_de_famille: Plagnol
    nom: Henri Plagnol
    type: depute
  depute_2430:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 2430
    adresses:
      - 24 Rue Gambetta 33230 Coutras Téléphone : 05 57 69 46 62 Télécopie : 05 57 69 46 63 
      - Permanence parlementaire 38 Bis Avenue de la République 33820 Braud-Saint-Louis Téléphone : 05 57 32 92 25 Télécopie : 05 57 64 53 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (11ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Plisson
    place_hemicycle: 643
    autresmandats:
      - Président de la Communauté de communes de l'Estuaire
      - Membre du conseil général (Gironde)
      - Maire de Saint-Caprais-de-Blaye, Gironde (405 habitants)
    mails:
      - philippe.plisson@free.fr
      - pplisson@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2430.asp
    profession: Retraité de l'enseignement
    site_web: http://www.philippeplisson.net
    debut_mandat: 20/06/2007
    nom: Philippe Plisson
    type: depute
  depute_2438:
    place_hemicycle: 262
    fonctions:
      - commission des affaires économiques / vice-président / 
    sexe: H
    id_an: 2438
    extras:
      - conseil de modération et de prévention / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2438.asp
    mails:
      - spoignant@assemblee-nationale.fr
      - serge.poignant@wanadoo.fr
    adresses:
      - Permanence parlementaire 290 Route du Loroux-Bottereau BP 22604 44115 Basse-Goulaine Téléphone : 02 40 06 20 57 Télécopie : 02 40 06 05 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Retraité du C.N.R.S.
    debut_mandat: 20/06/2007
    nom_de_famille: Poignant
    nom: Serge Poignant
    type: depute
  depute_243:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 243
    adresses:
      - Hôtel de ville 77410 Claye-Souilly Téléphone : 01 60 26 92 00 Télécopie : 01 60 26 30 06 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-et-Marne (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Albarello
    place_hemicycle: 225
    autresmandats:
      - Maire de Claye-Souilly, Seine-et-Marne (10152 habitants)
    mails:
      - yves.albarello@gmail.com
      - yalbarello@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/243.asp
    profession: Directeur administratif et financier
    site_web: http://www.albarello.info
    debut_mandat: 20/06/2007
    nom: Yves Albarello
    type: depute
  depute_2463:
    place_hemicycle: 111
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 2463
    mails:
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2463.asp
    circonscription: Pyrénées-Atlantiques (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur de société
    debut_mandat: 20/07/2007
    nom_de_famille: Poulou
    nom: Daniel Poulou
    type: depute
  depute_2473:
    fonctions:
      - commission des affaires sociales / vice-président / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 2473
    extras:
      - conseil de surveillance de la caisse nationale de l'assurance maladie des travailleurs salariés / membre titulaire
      - conseil de surveillance de la caisse nationale d'assurance vieillesse des travailleurs salariés / membre titulaire
      - conseil d'orientation des retraites / membre titulaire
    adresses:
      - 3 Place Napoléon 85000 La Roche-sur-Yon Téléphone : 02 51 37 87 70 Télécopie : 02 51 62 74 34 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vendée (1ère)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Préel
    place_hemicycle: 398
    mails:
      - jlpreel@orange.fr
      - jlpreel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2473.asp
    profession: Chef de service hospitalier
    site_web: http://www.preel.net
    debut_mandat: 20/06/2007
    nom: Jean-Luc Préel
    type: depute
  depute_2480:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2480
    extras:
      - conseil national pour le développement, l'aménagement et la protection de la montagne / membre titulaire
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Les Granges 43590 Beauzac Téléphone : 04 71 61 47 04 Télécopie : 04 71 61 47 10 
      - Permanence 2 Rue des Tanneries,  43000 Le Puy Téléphone : 04 71 02 16 44 Télécopie : 04 71 02 42 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 76 68 Télécopie : 01 40 63 79 66 
    circonscription: Haute-Loire (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Proriol
    place_hemicycle: 331
    autresmandats:
      - Maire de Beauzac, Haute-Loire (2493 habitants)
      - Membre du conseil régional (Auvergne)
    mails:
      - jproriol@assemblee-nationale.fr
      - mairie@ville-beauzac.fr
      - jproriol.permanence@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2480.asp
    profession: Ancien cadre
    site_web: http://www.bluebox.fr/jean-proriol
    debut_mandat: 20/06/2007
    nom: Jean Proriol
    type: depute
  depute_2492:
    fonctions:
      - commission des affaires européennes / vice-président / 
      - commission des lois / membre / 
    sexe: H
    id_an: 2492
    extras:
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre titulaire
    adresses:
      - 72 Avenue Charles de Gaulle 17620 Saint-Agnant Téléphone : 05 46 83 29 31 Télécopie : 05 46 39 11 15 
      - Permanence 21 Boulevard Germaine de la Falaise 17200 Royan Téléphone : 05 46 23 99 77 Télécopie : 05 46 39 11 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Charente-Maritime (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Quentin
    place_hemicycle: 267
    autresmandats:
      - Maire de Royan, Charente-Maritime (17102 habitants)
    mails:
      - dquentin@assemblee-nationale.fr
      - didierquentin@voila.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2492.asp
    profession: Ministre plénipotentiaire
    site_web: http://www.didierquentin.com
    debut_mandat: 20/06/2007
    nom: Didier Quentin
    type: depute
  depute_2494:
    place_hemicycle: 504
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Président du conseil régional (Rhône-Alpes)
    sexe: H
    id_an: 2494
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2494.asp
    mails:
      - jjqueyranne@assemblee-nationale.fr
    adresses:
      - 1 Rue Roger Salengro 69500 Bron Téléphone : 04 72 37 50 99 Télécopie : 04 72 37 58 87 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Maître de conférences à l'Université
    debut_mandat: 20/06/2007
    nom_de_famille: Queyranne
    nom: Jean-Jack Queyranne
    type: depute
  depute_2503:
    place_hemicycle: 480
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2503
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2503.asp
    mails:
      - dominiqueraimbourg@orange.fr
      - draimbourg@assemblee-nationale.fr
    adresses:
      - 73 Rue de la Commune de 1871 44400 Rezé  Téléphone : 02 40 02 73 80 Télécopie : 02 40 04 10 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Raimbourg
    nom: Dominique Raimbourg
    type: depute
  depute_2511:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2511
    adresses:
      - Mairie 121 Avenue de la Résistance 93340 Le Raincy Téléphone : 01 43 02 52 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Raoult
    place_hemicycle: 268
    autresmandats:
      - Maire du Raincy, Seine-Saint-Denis (12951 habitants)
    mails:
      - eraoult@assemblee-nationale.fr
      - ericraoult2007@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2511.asp
    profession: Assistant parlementaire du groupe RPR
    site_web: http://ericraoult.over-blog.com
    debut_mandat: 20/06/2007
    nom: Éric Raoult
    type: depute
  depute_2529:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2529
    adresses:
      - Mairie d'Altkirch 5 Place de la République 68130 Altkirch Téléphone : 03 89 40 00 04 Télécopie : 03 89 08 81 71 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 6 Place de la République 68130 Altkirch Téléphone : 03 89 40 17 75 Télécopie : 03 89 40 20 73 
    circonscription: Haut-Rhin (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Reitzer
    place_hemicycle: 166
    autresmandats:
      - Maire d'Altkirch, Haut-Rhin (5384 habitants)
    mails:
      - reitzer.jeanluc@free.fr
      - jlr.depute@online.fr
      - jlreitzer@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2529.asp
    profession: Cadre d'entreprise chargé des relations sociales
    site_web: http://www.depute-reitzer.net
    debut_mandat: 20/06/2007
    nom: Jean-Luc Reitzer
    type: depute
  depute_253:
    place_hemicycle: 123
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / membre / 
      - mission d'information commune sur les prix des carburants dans les dom / vice-président / 
    autresmandats:
      - Membre du Conseil municipal de Schoelcher, Martinique (20845 habitants)
    sexe: H
    id_an: 253
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/253.asp
    mails:
      - aalmont@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Martinique (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chargé de mission à la Chambre de Commerce et d'Industrie de la Martinique
    debut_mandat: 20/06/2007
    nom_de_famille: Almont
    nom: Alfred Almont
    type: depute
  depute_2549:
    place_hemicycle: 481
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 2549
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2549.asp
    mails:
      - mlreynaud@assemblee-nationale.fr
    adresses:
      - 44  Grand rue BP 40 16200 Jarnac Téléphone : 05 45 36 12 85 Télécopie : 05 45 82 28 81 
      - Téléphone mobile : 06 31 26 88 29  marie-line.reynaud@wanadoo.fr
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 69 88 (Téléphone assistant parlementaire) Téléphone : 01 40 63 69 74 Télécopie : 01 40 63 91 19  
    circonscription: Charente (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://marie-line-reynaud.parti-socialiste.fr/
    profession: Conseillère technique au centre d'information des droits de la femme
    debut_mandat: 20/06/2007
    nom_de_famille: Reynaud
    nom: Marie-Line Reynaud
    type: depute
  depute_2580:
    place_hemicycle: 80
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Adjoint au Maire de Marseille, Bouches-du-Rhône (798021 habitants)
    sexe: H
    id_an: 2580
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2580.asp
    mails:
      - jroatta@assemblee-nationale.fr
    adresses:
      - Mairie de Marseille 58 Boulevard Charles Livon Palais du Pharo 13007 Marseille Téléphone : 04 91 14 51 37 Télécopie : 04 91 14 51 67 
      - Permanence parlementaire 1 Rue de Suez 13007 Marseille Téléphone : 04 91 52 87 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Roatta
    nom: Jean Roatta
    type: depute
  depute_2591:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 2591
    extras:
      - conseil national pour le développement, l'aménagement et la protection de la montagne / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Résidence Destenay 3 Passage Bruzaud-Grille 65000 Tarbes Téléphone : 05 62 56 32 32 Télécopie : 05 62 34 83 65 
    circonscription: Hautes-Pyrénées (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Robin-Rodrigo
    place_hemicycle: 618
    autresmandats:
      - Vice-présidente du conseil général (Hautes-Pyrénées)
    mails:
      - c.robin-rodrigo@wanadoo.fr
      - crobin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2591.asp
    profession: Directeur départemental crédit immobilier
    site_web: http://chantalrobinrodrigo.hautetfort.com
    debut_mandat: 20/06/2007
    nom: Chantal Robin-Rodrigo
    type: depute
  depute_2597:
    fonctions:
      - commission des affaires étrangères / vice-président / 
    sexe: H
    id_an: 2597
    extras:
      - commission nationale pour l'élimination des mines antipersonnel / membre titulaire
      - conseil d'administration de l'agence pour l'enseignement français à l'étranger / membre titulaire
    adresses:
      - Permanence 4 Place Dorian BP 203 42408 Saint-Chamond cedex Téléphone : 04 77 31 46 55 Télécopie : 04 77 31 43 35 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (3ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Rochebloine
    place_hemicycle: 368
    autresmandats:
      - Vice-président du conseil général (Loire)
    mails:
      - frochebloine@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2597.asp
    profession: Directeur commercial
    site_web: http://www.francois-rochebloine.com
    debut_mandat: 20/06/2007
    nom: François Rochebloine
    type: depute
  depute_259:
    place_hemicycle: 87
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Vice-présidente du conseil régional (Basse Normandie)
    sexe: F
    id_an: 259
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/259.asp
    mails:
      - nameline@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire BP 20096 14603 Honfleur cedex Téléphone : 02 31 89 90 06 Télécopie : 02 31 89 32 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur territorial
    debut_mandat: 20/06/2007
    nom_de_famille: Ameline
    nom: Nicole Ameline
    type: depute
  depute_2600:
    fonctions:
      - commission des finances / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
    sexe: H
    id_an: 2600
    extras:
      - comité consultatif du secteur financier / membre suppléant
    adresses:
      - Hôtel de Ville 87031 Limoges cedex Téléphone : 05 55 45 60 00 Télécopie : 05 55 45 64 50 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Vienne (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Rodet
    place_hemicycle: 609
    autresmandats:
      - Maire de Limoges, Haute-Vienne (133907 habitants)
    mails:
      - arodet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2600.asp
    profession: Économiste
    debut_mandat: 20/06/2007
    nom: Alain Rodet
    type: depute
  depute_2603:
    fonctions:
      - commission des affaires culturelles et de l'éducation / vice-président / 
      - comité d'évaluation et de contrôle des politiques publiques / secrétaire / 
    sexe: H
    id_an: 2603
    adresses:
      - Permanence en circonscription 13 Boulevard Maréchal de Lattre de Tassigny 35000 Rennes Téléphone : 02 99 78 23 23 Télécopie : 02 99 59 78 02 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ille-et-Vilaine (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Rogemont
    place_hemicycle: 479
    autresmandats:
      - Membre du conseil général (Ille-et-Vilaine)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2603.asp
    mails:
      - marcel.rogemont@wanadoo.fr
    site_web: http://www.marcelrogemont.net
    profession: Cadre
    debut_mandat: 20/06/2007
    nom: Marcel Rogemont
    type: depute
  depute_2608:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 2608
    adresses:
      - Mairie 84045 Avignon cedex Téléphone : 04 90 80 83 85 Télécopie : 04 90 80 83 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vaucluse (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Roig
    place_hemicycle: 192
    autresmandats:
      - Maire d'Avignon, Vaucluse (85929 habitants)
    mails:
      - mjroig@assemblee-nationale.fr
      - marie-josee.roig@mairie-avignon.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2608.asp
    profession: Professeur de lettres
    site_web: http://www.mjroig.fr
    debut_mandat: 20/06/2007
    nom: Marie-Josée Roig
    type: depute
  depute_2611:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2611
    adresses:
      - Permanence 165 Rue d'Arras 59000 Lille Téléphone : 03 20 52 09 20 Télécopie : 03 28 54 01 37 
      - Conseil régional Hôtel de Région, Centre Rihour 59555 Lille cedex 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Roman
    place_hemicycle: 510
    autresmandats:
      - Vice-président du conseil régional (Nord-Pas-de-Calais)
    mails:
      - contact@bernard-roman.org
      - broman@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2611.asp
    profession: Avocat, administrateur territorial
    site_web: http://www.bernard-roman.net
    debut_mandat: 20/06/2007
    nom: Bernard Roman
    type: depute
  depute_2631:
    place_hemicycle: 467
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Vice-président de la communauté d'agglomération de la plaine centrale du Val-de-Marne
      - Maire d'Alfortville, Val-de-Marne (36151 habitants)
    sexe: H
    id_an: 2631
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2631.asp
    mails:
      - rrouquet@assemblee-nationale.fr
    adresses:
      - Mairie 94140 Alfortville Téléphone : 01 58 73 29 00 Télécopie : 01 43 75 07 64 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (9ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Électromécanicien
    debut_mandat: 20/06/2007
    nom_de_famille: Rouquet
    nom: René Rouquet
    type: depute
  depute_2640:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 2640
    adresses:
      - Permanence parlementaire 8 Rue Jules Cazot 30100 Alès  Téléphone : 04 66 52 01 89 Télécopie : 04 66 52 01 13 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gard (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Roustan
    place_hemicycle: 140
    autresmandats:
      - Maire d'Alès, Gard (39346 habitants)
      - Président de la Communauté d'Agglomération du Grand Alès en Cévennes
    mails:
      - mroustan@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2640.asp
    profession: Professeur d'enseignement technique
    site_web: http://maxroustan.fr
    debut_mandat: 20/06/2007
    nom: Max Roustan
    type: depute
  depute_265:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 265
    adresses:
      - Permanence  28 Avenue Charles de Gaulle 71400 Autun Téléphone : 03 85 52 31 45 Télécopie : 03 85 86 10 46 
      - Permanence 14 Rue du Maréchal Leclerc 71200 Le Creusot Téléphone : 03 85 55 60 47 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Anciaux
    place_hemicycle: 195
    autresmandats:
      - Membre du Conseil municipal d'Autun, Saône-et-Loire (16432 habitants)
      - Membre du conseil régional (Bourgogne)
    mails:
      - jpanciaux@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/265.asp
    profession: Technicien qualiticien
    site_web: http://www.jeanpaulanciaux.com
    debut_mandat: 20/06/2007
    nom: Jean-Paul Anciaux
    type: depute
  depute_2661:
    place_hemicycle: 518
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Mérignac, Gironde (61992 habitants)
      - Vice-président de la communauté urbaine de Bordeaux
    sexe: H
    id_an: 2661
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2661.asp
    mails:
      - msainte@assemblee-nationale.fr
    adresses:
      - Boîte postale 20154 33706 Mérignac cedex Téléphone : 05 56 55 66 15 Téléphone : 05 56 55 66 10 Télécopie : 05 56 55 66 06 Télécopie : 05 56 55 66 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Sainte-Marie
    nom: Michel Sainte-Marie
    type: depute
  depute_266776:
    place_hemicycle: 216
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Maire de Niederbronn-les-Bains, Bas-Rhin (4319 habitants)
    sexe: H
    id_an: 266776
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266776.asp
    mails:
      - freiss@assemblee-nationale.fr
      - reiss.depute@wanadoo.fr
    adresses:
      - Permanence parlementaire 12 Allée des Peupliers BP 2 67161 Wissembourg cedex Téléphone : 03 88 54 81 00 Télécopie : 03 88 94 18 16 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Agrégé de mathématiques
    debut_mandat: 20/06/2007
    nom_de_famille: Reiss
    nom: Frédéric Reiss
    type: depute
  depute_266782:
    place_hemicycle: 20
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Sablé-sur-Sarthe, Sarthe (12716 habitants)
      - Vice-président de la communauté de communes du district de Sablé sur Sarthe
    sexe: H
    id_an: 266782
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266782.asp
    circonscription: Sarthe (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/07/2007
    nom_de_famille: Joulaud
    nom: Marc Joulaud
    type: depute
  depute_266788:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / membre / 
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission des lois / membre / 
    sexe: H
    id_an: 266788
    extras:
      - comité de surveillance de l'établissement de gestion du fonds de financement des prestations sociales des non-salariés agricoles / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 35 Télécopie :  01 40 63 32 84 
      - Hôtel de la paix Avenue Brazza 48100 Marvejols Téléphone : 04 66 32 08 09 Télécopie : 04 66 32 08 10 
      - Mairie 48310 Fournels Téléphone : 04 66 31 60 15 Télécopie : 04 66 31 60 13 
    circonscription: Lozère (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Morel-A-L'Huissier
    place_hemicycle: 137
    autresmandats:
      - Membre du conseil général (Lozère)
      - Président de la communauté de communes des Hautes Terres
      - Maire de Fournels, Lozère (324 habitants)
    mails:
      - pmorelalhuissier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266788.asp
    profession: Avocat
    site_web: http://www.pierre-morel.fr
    debut_mandat: 20/06/2007
    nom: Pierre Morel-A-L'Huissier
    type: depute
  depute_266793:
    place_hemicycle: 17
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Vice-président du conseil général (Cantal)
      - Maire d'Ally, Cantal (701 habitants)
    sexe: H
    id_an: 266793
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266793.asp
    circonscription: Cantal (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Exploitant agricole
    debut_mandat: 20/07/2007
    nom_de_famille: Bony
    nom: Jean-Yves Bony
    type: depute
  depute_266797:
    fonctions:
      - commission des lois / secrétaire / 
    sexe: H
    id_an: 266797
    extras:
      - commission supérieure de codification / membre titulaire
      - commission nationale de l'informatique et des libertés / membre titulaire
    adresses:
      - Permanence parlementaire 45 Route de Villedieu 50000 Saint Lô Téléphone : 02 33 05 05 50 Télécopie : 02 33 57 39 98 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Manche (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gosselin
    place_hemicycle: 150
    autresmandats:
      - Président de la communauté de communes de Marigny
      - Maire de Remilly-sur-Lozon, Manche (556 habitants)
    mails:
      - pgosselin@assemblee-nationale.fr
      - philippegosselin50@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266797.asp
    profession: Professeur de droit en classes préparatoires aux grandes écoles
    site_web: http://www.philippegosselin.fr
    debut_mandat: 20/06/2007
    nom: Philippe Gosselin
    type: depute
  depute_2667:
    fonctions:
      - assemblée nationale / vice-président / 27/06/2007
      - délégation chargée de la communication et de la presse / membre / 
      - délégation chargée de l'informatique et des nouvelles technologies / président / 
      - délégation chargée des activités internationales / membre / 
      - délégation chargée des représentants d'intérêts / membre / 
      - commission des affaires étrangères / membre / 
      - délégation spéciale chargée de la question des groupes d'intérêt / membre / 
      - délégation chargée de l'application du statut du député / membre / 
      - délégation chargée de la communication audiovisuelle et de la presse / membre / 
    sexe: H
    id_an: 2667
    adresses:
      - 31 Avenue Jean Médecin 06000 Nice Téléphone : 04 93 80 35 00 Télécopie : 04 93 80 02 56 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-Maritimes (3ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Salles
    place_hemicycle: 365
    autresmandats:
      - Membre du conseil régional (Provence-Alpes-Côte-d'Azur)
      - Adjoint au Maire de Nice, Alpes-Maritimes (342482 habitants)
    mails:
      - contact@rudy-salles.com
      - rsalles@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2667.asp
    profession: Avocat
    site_web: http://www.rudy-salles.com
    debut_mandat: 20/06/2007
    nom: Rudy Salles
    type: depute
  depute_266815:
    fonctions:
      - commission des affaires économiques / membre / 
      - mission d'information commune sur les prix des carburants dans les dom / rapporteur / 
    sexe: H
    id_an: 266815
    extras:
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre suppléant
      - conseil national du littoral / membre titulaire
    adresses:
      - Permanence 54 Quai de Léon 29800 Landerneau Téléphone : 02 98 85 66 96 Télécopie : 02 98 21 58 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Finistère (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Guen
    place_hemicycle: 120
    autresmandats:
      - Membre du conseil général (Finistère)
      - Président de la communauté de communes de la Baie du Kernic
      - Membre du Conseil municipal de Plounévez-Lochrist, Finistère (2278 habitants)
    mails:
      - jleguen@assemblee-nationale.fr
      - jacques-leguen@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/266815.asp
    profession: Docteur en médecine
    site_web: http://www.jacquesleguen.org
    debut_mandat: 20/06/2007
    nom: Jacques Le Guen
    type: depute
  depute_267003:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267003
    extras:
      - haut conseil du secteur public / membre titulaire
      - conseil supérieur des prestations sociales agricoles / membre suppléant
    adresses:
      - Rue de Salassous 48700 Rieutort-de-Randon Téléphone : 04 66 47 19 79 
      - 1 Rue des Carces 48000 Mende 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Lozère (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Saint-Léger
    place_hemicycle: 227
    autresmandats:
      - Membre du conseil régional (Languedoc-Roussillon)
    mails:
      - contact@francissaintleger.fr
      - fsaint@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267003.asp
    profession: Ingénieur
    debut_mandat: 20/06/2007
    nom: Francis Saint-Léger
    type: depute
  depute_267013:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267013
    adresses:
      - Permanence parlementaire 3 Faubourg de Belfort 68700 Cernay Téléphone : 03 89 75 83 95 Télécopie : 03 89 75 63 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Sordi
    place_hemicycle: 301
    autresmandats:
      - Président de la communauté de communes de Cernay-et-Environs
      - Maire de Cernay, Haut-Rhin (10446 habitants)
    mails:
      - michel.sordi.depute@wanadoo.fr
      - msordi@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267013.asp
    profession: Cadre d'entreprise
    site_web: http://michel.sordi.over-blog.com
    debut_mandat: 20/06/2007
    nom: Michel Sordi
    type: depute
  depute_267018:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / secrétaire / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267018
    extras:
      - conseil supérieur des prestations sociales agricoles / membre titulaire
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Permanence parlementaire 13  Rue de la Tour BP 50056 70302 Luxeuil-les-Bains cedex Téléphone : 03 84 40 62 35 Télécopie : 03 84 40 35 05 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Saône (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Raison
    place_hemicycle: 2
    autresmandats:
      - Maire de Luxeuil-les-Bains, Haute-Saône (8416 habitants)
    mails:
      - michel.raison@michel-raison.net
      - mraison@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267018.asp
    profession: Agriculteur
    site_web: http://www.michelraison.fr
    debut_mandat: 20/06/2007
    nom: Michel Raison
    type: depute
  depute_267028:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267028
    adresses:
      - Permanence  21 Rue des Mégissiers BP 21 76290 Montivilliers Téléphone : 02 35 20 74 55 Télécopie : 02 35 55 28 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 28 Rue de l'Inondation BP 61 76400 Fécamp Téléphone : 02 35 28 53 09 Télécopie : 02 35 27 79 86 
    circonscription: Seine-Maritime (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Fidelin
    place_hemicycle: 141
    autresmandats:
      - Maire de Mannevillette, Seine-Maritime (690 habitants)
      - Vice-président de la communauté de l'Agglomération Havraise
      - Membre du conseil général (Seine-Maritime)
    mails:
      - dfidelin@assemblee-nationale.fr
      - fidelin.monti@wanadoo.fr
      - d.fidelin.depute@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267028.asp
    profession: Assureur
    site_web: http://www.danielfidelin.net
    debut_mandat: 20/06/2007
    nom: Daniel Fidelin
    type: depute
  depute_267031:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267031
    extras:
      - conseil supérieur de l'énergie / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 14 Rue Albert Bochet 76440 Forges-les-Eaux Téléphone : 02 35 09 36 53 Télécopie : 02 35 09 36 57 
    circonscription: Seine-Maritime (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lejeune
    place_hemicycle: 211
    autresmandats:
      - Maire de Forges-les-Eaux, Seine-Maritime (3461 habitants)
      - Membre du conseil général (Seine-Maritime)
    mails:
      - mlejeune@assemblee-nationale.fr
      - mlejeune.depute76@wanadoo.fr
      - mlejeune@forgesleseaux.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267031.asp
    profession: Vétérinaire
    debut_mandat: 20/06/2007
    nom: Michel Lejeune
    type: depute
  depute_267042:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267042
    adresses:
      - 6 Boulevard du Général Leclerc 53100 Mayenne Téléphone : 02 43 30 29 60 Télécopie : 02 43 30 29 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Mayenne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Favennec
    place_hemicycle: 339
    autresmandats:
      - Membre du conseil régional (Pays de la Loire)
    mails:
      - yfavennec@assemblee-nationale.fr
      - favennec.yannick@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267042.asp
    profession: Directeur de cabinet
    site_web: http://www.yannickfavennec.com
    debut_mandat: 20/06/2007
    nom: Yannick Favennec
    type: depute
  depute_267049:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267049
    adresses:
      - Permanence parlementaire 3 Allée Forestière BP 40122 56501 Locminé cedex Téléphone : 02 97 60 09 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Morbihan (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lorgeoux
    place_hemicycle: 32
    autresmandats:
      - Vice-président du conseil général (Morbihan)
    mails:
      - glorgeoux@assemblee-nationale.fr
      - gerardlorgeouxdepute@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267049.asp
    profession: Imprimeur
    site_web: http://www.gerardlorgeoux.com
    debut_mandat: 20/06/2007
    nom: Gérard Lorgeoux
    type: depute
  depute_267057:
    place_hemicycle: 222
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire de Sarreguemines, Moselle (23202 habitants)
    sexe: H
    id_an: 267057
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267057.asp
    mails:
      - clett@assemblee-nationale.fr
      - clett@wanadoo.fr
    adresses:
      - Permanence 18A Rue Chamborand 57200 Sarreguemines Téléphone : 03 87 98 33 68 Télécopie : 03 87 98 36 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Moselle (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre hospitalier
    debut_mandat: 20/06/2007
    nom_de_famille: Lett
    nom: Céleste Lett
    type: depute
  depute_267069:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / vice-président / 
      - comité d'évaluation et de contrôle des politiques publiques / vice-président / 
      - mission d'information commune sur les exonérations sociales / membre / 
    sexe: H
    id_an: 267069
    extras:
      - conseil national de l'aménagement et du développement du territoire / membre titulaire
      - comité consultatif de la législation et de la réglementation financières / membre titulaire
      - conseil d'administration de l'établissement public "autoroutes de france" / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 29 Boulevard Berthelot 63400 Chamalières Téléphone : 04 73 19 19 73 Télécopie : 04 73 36 24 16 
    circonscription: Puy-de-Dôme (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: d'Estaing
    place_hemicycle: 286
    autresmandats:
      - Maire de Chamalières, Puy-de-Dôme (18134 habitants)
    mails:
      - louis.giscard-destaing@wanadoo.fr
      - lgiscarddestaing@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267069.asp
    profession: Chef d'entreprise
    site_web: http://www.lge-pour-clermontmontagne.fr
    debut_mandat: 20/06/2007
    nom: Louis Giscard d'Estaing
    type: depute
  depute_267075:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 267075
    extras:
      - commission supérieure de codification / membre suppléant
      - conseil d'orientation de la simplification administrative / membre titulaire
    adresses:
      - Mairie 73 Avenue des Thermes 01220 Divonne-les-Bains Téléphone : 04 50 99 17 45 Télécopie : 04 50 99 16 75 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ain (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Blanc
    place_hemicycle: 45
    autresmandats:
      - Président de la communauté de communes du Pays de Gex
      - Maire de Divonne-les-Bains, Ain (6171 habitants)
    mails:
      - contact@etienne-blanc.org
      - eblanc@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267075.asp
    profession: Avocat
    site_web: http://www.etienne-blanc.org
    debut_mandat: 20/06/2007
    nom: Étienne Blanc
    type: depute
  depute_267080:
    place_hemicycle: 88
    fonctions:
      - commission des finances / membre / 
      - mandat de député suite à la cessation de fonction de membre du gouvernement le : 15/02/2009 / reprise de l'exercice / 
    autresmandats:
      - Membre de la Communauté d'agglomération de Saint-Quentin
      - Adjoint au Maire de Saint-Quentin, Aisne (59066 habitants)
    sexe: H
    id_an: 267080
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267080.asp
    mails:
      - xbertrand@assemblee-nationale.fr
    adresses:
      - Permanence 19 Rue du Gouvernement 02100 Saint-Quentin Téléphone : 03 23 05 22 66 Télécopie : 03 23 05 41 74 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aisne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Agent d'assurance
    debut_mandat: 20/06/2007
    nom_de_famille: Bertrand
    nom: Xavier Bertrand
    type: depute
  depute_267087:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / vice-président / 
    sexe: H
    id_an: 267087
    extras:
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Permanence parlementaire 2 Rue Pierre Courbet 47000 Agen Téléphone : 05 53 67 87 61 Télécopie : 05 53 95 58 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 71 76 Téléphone : 06 19 89 00 32 Télécopie : 01 40 63 78 04 
    circonscription: Lot-et-Garonne (1ère)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Séjour
    place_hemicycle: 397
    autresmandats:
      - Président de la Communauté d'agglomération d'Agen
      - Maire d'Agen, Lot-et-Garonne (30099 habitants)
    mails:
      - jdionisdusejour@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267087.asp
    profession: Ingénieur
    site_web: http://www.jeandionis.com
    debut_mandat: 20/06/2007
    nom: Jean Dionis du Séjour
    type: depute
  depute_267091:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 267091
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ariège (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Massat
    place_hemicycle: 569
    autresmandats:
      - Membre du Conseil municipal de Foix, Ariège (9109 habitants)
    mails:
      - fmassat@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267091.asp
    profession: Fonctionnaire territoriale
    site_web: http://www.frederiquemassat.com
    debut_mandat: 20/06/2007
    nom: Frédérique Massat
    type: depute
  depute_267099:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267099
    extras:
      - conseil supérieur de l'établissement national des invalides de la marine / membre titulaire
    adresses:
      - Villa Molière 19 Place Saint-Patrice BP 53501 14405 Bayeux cedex Téléphone : 02 31 51 73 73 Télécopie : 02 31 22 91 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lefranc
    place_hemicycle: 109
    autresmandats:
      - Membre du conseil régional (Basse Normandie)
    mails:
      - jmlefrancdepute@wanadoo.fr
      - jmlefranc@assemblee-nationale.fr
      - contact@jmlefranc.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267099.asp
    site_web: http://www.jmlefranc.fr
    debut_mandat: 20/06/2007
    nom: Jean-Marc Lefranc
    type: depute
  depute_267110:
    place_hemicycle: 389
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Membre du conseil général (Eure)
      - Maire de Beaumesnil, Eure (560 habitants)
    sexe: H
    id_an: 267110
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267110.asp
    circonscription: Eure (3ème)
    groupe:
      - nouveau centre / membre
    profession: Informaticien retraité
    debut_mandat: 20/07/2007
    nom_de_famille: Vampa
    nom: Marc Vampa
    type: depute
  depute_267118:
    fonctions:
      - commission de la défense nationale et des forces armées / secrétaire / 
    sexe: H
    id_an: 267118
    adresses:
      - 2 Rue Amiral Bauguen 29150 Châteaulin Téléphone : 02 98 86 66 20  Télécopie : 02 98 86 66 26 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Finistère (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ménard
    place_hemicycle: 51
    autresmandats:
      - Maire de Châteauneuf-du-Faou, Finistère (3595 habitants)
    mails:
      - cmenard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267118.asp
    profession: Médecin
    site_web: http://cmenard.com
    debut_mandat: 20/06/2007
    nom: Christian Ménard
    type: depute
  depute_267140:
    place_hemicycle: 14
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Membre du conseil général (Drôme)
      - Maire de Hauterives, Drôme (1333 habitants)
    sexe: H
    id_an: 267140
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267140.asp
    mails:
      - gabriel.biancheri@wanadoo.fr
      - gbiancheri@assemblee-nationale.fr
    adresses:
      - Permanence 23 Rue Jacquemart 26100 Romans Téléphone : 04 75 05 19 62 Télécopie : 04 75 05 19 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Drôme (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Vétérinaire
    debut_mandat: 20/06/2007
    nom_de_famille: Biancheri
    nom: Gabriel Biancheri
    type: depute
  depute_267144:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267144
    extras:
      - conseil supérieur de l'énergie / membre titulaire
    adresses:
      - Permanence 2 Rue de la Petite Cité BP 146 27001 Évreux cedex Téléphone : 02 32 38 74 07 Télécopie : 02 32 33 69 90 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Eure (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Nicolas
    place_hemicycle: 281
    autresmandats:
      - Membre du Conseil municipal d'Évreux, Eure (51226 habitants)
    mails:
      - jpnicolas@assemblee-nationale.fr
      - jean.pierre.nicolas@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267144.asp
    profession: Ingénieur
    site_web: http://www.jean-pierre-nicolas.fr
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Nicolas
    type: depute
  depute_267148:
    place_hemicycle: 133
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267148
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267148.asp
    mails:
      - fgilard@assemblee-nationale.fr
    adresses:
      - 1 Rue Turnèbe 27700 Les Andelys Téléphone : 02 32 64 20 95 Télécopie : 02 32 71 06 24 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Eure (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.franckgilard.info 
    profession: Consultant
    debut_mandat: 20/06/2007
    nom_de_famille: Gilard
    nom: Franck Gilard
    type: depute
  depute_267151:
    place_hemicycle: 340
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    autresmandats:
      - Président de la communauté d'agglomération "Chartres Métropole"
      - Maire de Chartres, Eure-et-Loir (40431 habitants)
    sexe: H
    id_an: 267151
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267151.asp
    circonscription: Eure-et-Loir (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur informatique
    debut_mandat: 15/09/2008
    nom_de_famille: Gorges
    nom: Jean-Pierre Gorges
    type: depute
  depute_267166:
    place_hemicycle: 380
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Première adjointe de Langres, Haute-Marne (9586 habitants)
    sexe: F
    id_an: 267166
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267166.asp
    circonscription: Haute-Marne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin du travail
    debut_mandat: 20/07/2007
    nom_de_famille: Delong
    nom: Sophie Delong
    type: depute
  depute_267178:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267178
    adresses:
      - 7 Rue Joseph Gaucher 10500 Brienne-le-Château Téléphone : 03 25 92 20 31 Télécopie : 03 25 92 22 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 19 43 Télécopie : 01 40 63 19 45 
      - Mairie Place de l'Hôtel de ville 10500 Brienne-le-Château Téléphone : 03 25 92 80 31 
    circonscription: Aube (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Dhuicq
    place_hemicycle: 239
    autresmandats:
      - Maire de Brienne le Château, Aube (3336 habitants)
      - Membre du conseil général (Aube)
    mails:
      - ndhuicq@orange.fr
      - ndhuicq@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267178.asp
    profession: Psychiatre des hôpitaux
    site_web: http://www.nicolasdhuicq.com
    debut_mandat: 20/06/2007
    nom: Nicolas Dhuicq
    type: depute
  depute_267182:
    place_hemicycle: 122
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Maire de Vire, Calvados (12815 habitants)
    sexe: H
    id_an: 267182
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267182.asp
    mails:
      - jycousin@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville 14500 Vire Téléphone : 02 31 68 99 47 Téléphone : 02 31 66 60 00 Télécopie : 02 31 67 37 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Inspecteur principal des impôts
    debut_mandat: 20/06/2007
    nom_de_famille: Cousin
    nom: Jean-Yves Cousin
    type: depute
  depute_267188:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 267188
    extras:
      - conseil de surveillance du fonds de financement de la protection complémentaire  de la couverture universelle du risque maladie / membre titulaire
      - conseil supérieur pour le reclassement professionnel et social des travailleurs handicapés / membre titulaire
    adresses:
      - 1 Bis Avenue Saint Just 58000 Nevers Téléphone : 03 86 61 80 90 Télécopie : 03 86 36 53 47 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville Place de l'Hôtel de Ville 58000 Nevers Téléphone : 03 86 68 46 03 
    circonscription: Nièvre (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Carrillon-Couvreur
    place_hemicycle: 361
    autresmandats:
      - Adjointe au Maire de Nevers, Nièvre (40932 habitants)
    mails:
      - mcarrillon@assemblee-nationale.fr
      - martine-carrillon@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267188.asp
    profession: Directrice d'un institut médico-éducatif
    debut_mandat: 20/06/2007
    nom: Martine Carrillon-Couvreur
    type: depute
  depute_2671:
    place_hemicycle: 587
    fonctions:
      - commission des finances / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - bureau du comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: H
    id_an: 2671
    extras:
      - conseil supérieur de la réserve militaire / membre suppléant
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2671.asp
    mails:
      - jcsandrier@assemblee-nationale.fr
      - JC.SANDRIER@wanadoo.fr
    adresses:
      - 7 Avenue de la République 18100 Vierzon Téléphone : 02 48 52 28 43 Télécopie : 02 48 52 28 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Cher (2ème)
    groupe:
      - gauche démocrate et républicaine / président
    profession: Chimiste
    debut_mandat: 20/06/2007
    nom_de_famille: Sandrier
    nom: Jean-Claude Sandrier
    type: depute
  depute_267200:
    fonctions:
      - commission des lois / secrétaire / 
    sexe: H
    id_an: 267200
    extras:
      - commission nationale de l'informatique et des libertés / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 234 Rue du Général de Gaulle 59139 Wattignies Téléphone : 03 20 60 26 26 Télécopie : 03 20 60 38 34 
    circonscription: Nord (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Huyghe
    place_hemicycle: 200
    autresmandats:
      - Membre de la communauté urbaine de Lille Métropole
      - Membre du Conseil municipal de Lille, Nord (184231 habitants)
    mails:
      - hr.huyghe@orange.fr
      - shuyghe@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267200.asp
    profession: Notaire
    site_web: http://sebastienhuyghe.blogs.com 
    debut_mandat: 20/06/2007
    nom: Sébastien Huyghe
    type: depute
  depute_267204:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267204
    adresses:
      - 39  Grande Rue 39600 Cramans Téléphone : 03 84 37 72 49 Télécopie : 03 84 37 68 40 
      - 17 Rue Marcel Aymé 39100 Dole Téléphone : 03 84 72 08 01 Télécopie : 03 84 82 07 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 32 67 Téléphone : 01 40 63 32 17 Télécopie : 01 40 63 32 97 
    circonscription: Jura (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Sermier
    place_hemicycle: 309
    autresmandats:
      - Maire de Cramans, Jura (429 habitants)
      - Membre du conseil général (Jura)
    mails:
      - jmsermier@assemblee-nationale.fr
      - jmsermier-dole@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267204.asp
    profession: Viticulteur
    site_web: http://jm-sermier.fr
    debut_mandat: 20/06/2007
    nom: Jean-Marie Sermier
    type: depute
  depute_267209:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 267209
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 01 56 Téléphone : 01 40 63 01 06 Télécopie : 01 40 63 01 86 
    circonscription: Loir-et-Cher (1ère)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Perruchot
    place_hemicycle: 374
    autresmandats:
      - Membre du Conseil municipal de Blois, Loir-et-Cher (49184 habitants)
    mails:
      - nperruchot@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267209.asp
    profession: Consultant en entreprise
    site_web: http://nicolasperruchot.fr/
    debut_mandat: 20/06/2007
    nom: Nicolas Perruchot
    type: depute
  depute_267224:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / vice-président / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267224
    adresses:
      - Hôtel de Ville Avenue Pablo Casals 66450 Pollestres Téléphone : 04 68 85 70 75 Télécopie : 04 68 85 70 77 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Orientales (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mach
    place_hemicycle: 147
    autresmandats:
      - Maire de Pollestres, Pyrénées-Orientales (3623 habitants)
      - Vice-président de la Communauté d'agglomération Perpignan Méditerranée
    mails:
      - dmach@assemblee-nationale.fr
      - daniel.mach@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267224.asp
    profession: Cadre commercial
    site_web: http://www.danielmach.fr
    debut_mandat: 20/06/2007
    nom: Daniel Mach
    type: depute
  depute_267227:
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - délégation chargée des représentants d'intérêts / membre / 
      - commission des finances / membre / 
      - délégation chargée de l'application du statut du député / membre / 
      - assemblée nationale / secrétaire / 01/10/2008
    sexe: F
    id_an: 267227
    extras:
      - conseil supérieur du service public ferroviaire / membre titulaire
      - commission de surveillance de la caisse des dépôts et consignations / membre titulaire
    adresses:
      - Permanence 26B Rue de la Wanne 68100 Mulhouse Téléphone : 03 89 31 70 00 Télécopie : 03 89 44 65 23 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Grosskost
    place_hemicycle: 282
    autresmandats:
      - Vice-présidente du conseil régional (Alsace)
    mails:
      - agrosskost@assemblee-nationale.fr
      - depute.grosskost@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267227.asp
    profession: Avocat
    site_web: http://www.arlette-grosskost.com
    debut_mandat: 20/06/2007
    nom: Arlette Grosskost
    type: depute
  depute_267233:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267233
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Place Jean Jaurès 76380 Canteleu Téléphone : 02 35 23 57 89 Télécopie : 02 35 36 44 70 
    circonscription: Seine-Maritime (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bouillon
    place_hemicycle: 634
    autresmandats:
      - Maire de Canteleu, Seine-Maritime (15429 habitants)
    mails:
      - cbouillon@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267233.asp
    profession: Fonctionnaire de catégorie A
    site_web: http://www.christophebouillon.fr
    debut_mandat: 20/06/2007
    nom: Christophe Bouillon
    type: depute
  depute_267241:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / vice-président / 
    sexe: H
    id_an: 267241
    extras:
      - conseil national du bruit / membre titulaire
    adresses:
      - Hôtel de Ville, Cabinet du Maire Place Émile Leturcq 80300 Albert Téléphone : 03 22 74 38 51 Télécopie : 03 22 74 38 58 
      - Permanence parlementaire Rue de la Caisse d'épargne 80200 Péronne Téléphone : 03 22 84 38 43 Télécopie : 03 22 84 37 43 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Somme (5ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Demilly
    place_hemicycle: 386
    autresmandats:
      - Président de la communauté de communes du Pays du Coquelicot
      - Maire d'Albert, Somme (10065 habitants)
    mails:
      - depute.demilly@wanadoo.fr
      - sdemilly@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267241.asp
    profession: Consultant en management
    site_web: http://www.stephane-demilly.org
    debut_mandat: 20/06/2007
    nom: Stéphane Demilly
    type: depute
  depute_267246:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267246
    adresses:
      - Permanence parlementaire 11 Rue de la Préfecture 88000 Épinal Téléphone : 03 29 35 76 25 Télécopie : 03 29 82 95 57 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie Rue du Général Leclerc 88000 Épinal Téléphone : 03 29 68 50 15 Télécopie : 03 29 34 16 06 
    circonscription: Vosges (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Heinrich
    place_hemicycle: 118
    autresmandats:
      - Maire d'Épinal, Vosges (35788 habitants)
    mails:
      - mheinrich@assemblee-nationale.fr
      - michelheinrich.depute@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267246.asp
    profession: Pharmacien
    site_web: http://www.michel-heinrich.fr
    debut_mandat: 20/06/2007
    nom: Michel Heinrich
    type: depute
  depute_267253:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267253
    adresses:
      - 8 Place Saint-Pierre 04400 Barcelonnette Téléphone : 04 92 81 42 45 
      - Mairie 04200 Sisteron Téléphone : 04 92 61 40 71 Télécopie : 04 92 61 56 59 
      - 171  Avenue Paul Arène BP 25 04201 Sisteron cedex 01 Téléphone : 04 92 61 40 71 Télécopie : 04 92 61 56 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-de-Haute-Provence (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Spagnou
    place_hemicycle: 116
    autresmandats:
      - Maire de Sisteron, Alpes-de-Haute-Provence (6964 habitants)
      - Président de la communauté de communes du Sisteronais
    mails:
      - dspagnou@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267253.asp
    profession: Directeur de caisse d'épargne retraité
    site_web: http://www.danielspagnou.com
    debut_mandat: 20/06/2007
    nom: Daniel Spagnou
    type: depute
  depute_267257:
    place_hemicycle: 293
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Maire de Vals-les-Bains, Ardèche (3536 habitants)
    sexe: H
    id_an: 267257
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267257.asp
    mails:
      - jcflory@assemblee-nationale.fr
      - jean-claude.flory@wanadoo.fr
    adresses:
      - Permanence parlementaire BP 107 07600 Vals les Bains Téléphone : 04 75 37 90 25 Télécopie : 04 75 38 07 16 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ardèche (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Conseiller en gestion locale
    debut_mandat: 20/06/2007
    nom_de_famille: Flory
    nom: Jean-Claude Flory
    type: depute
  depute_267260:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / secrétaire / 
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 267260
    extras:
      - conseil de surveillance du fonds de réserve pour les retraites / membre suppléante
      - commision nationale d'agrément des associations représentant les usagers dans les instances hospitalières ou de santé publique / membre titulaire
    adresses:
      - Permanence parlementaire 21 Avenue du Maréchal Leclerc 08000 Charleville-Mézières Téléphone : 03 24 32 49 81 Télécopie : 03 24 33 92 16 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ardennes (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Poletti
    place_hemicycle: 92
    autresmandats:
      - Membre du conseil régional (Champagne-Ardenne)
    mails:
      - bpoletti@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267260.asp
    profession: Sage-femme
    site_web: http://www.berengere-poletti.fr
    debut_mandat: 20/06/2007
    nom: Bérengère Poletti
    type: depute
  depute_267266:
    fonctions:
      - commission des finances / vice-président / 
    sexe: H
    id_an: 267266
    extras:
      - conseil supérieur des prestations sociales agricoles / membre suppléant
      - conseil national de l'enseignement supérieur privé / membre suppléant
    adresses:
      - 5 Boulevard de la République 12000 Rodez Téléphone : 05 65 67 51 00 Télécopie : 05 65 67 00 44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aveyron (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Censi
    place_hemicycle: 79
    mails:
      - ycensi@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267266.asp
    profession: Ingénieur conseil
    site_web: http://www.yvescensi.com
    debut_mandat: 20/06/2007
    nom: Yves Censi
    type: depute
  depute_267270:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 267270
    extras:
      - comité national d'évaluation des dispositifs expérimentaux d'aide aux personnes âgées / membre suppléant
      - comité national de l'organisation sanitaire et sociale / membre suppléant
    adresses:
      - Hôtel de Ville Place Guillaume-le-Conquérant 14700 Falaise Téléphone : 02 31 41 66 85 Télécopie : 02 31 20 02 92 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Calvados (3ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Leteurtre
    place_hemicycle: 401
    autresmandats:
      - Vice-président du conseil général (Calvados)
    mails:
      - cleteurtre@falaise.fr
      - cleteurtre@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267270.asp
    profession: Chirurgien orthopédiste
    site_web: http://www.claudeleteurtre.net
    debut_mandat: 20/06/2007
    nom: Claude Leteurtre
    type: depute
  depute_267278:
    place_hemicycle: 517
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Président du conseil général (Gers)
    sexe: H
    id_an: 267278
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267278.asp
    mails:
      - pmartin@cg32.fr
      - pmartin@assemblee-nationale.fr
      - ph.martin-depute@wanadoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 81  Route de Pessan 32000 Auch Téléphone : 05 62 63 44 48 Télécopie : 05 62 63 46 85 
    circonscription: Gers (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Préfet
    debut_mandat: 20/06/2007
    nom_de_famille: Martin
    nom: Philippe Martin
    type: depute
  depute_267283:
    place_hemicycle: 59
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267283
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267283.asp
    circonscription: Indre-et-Loire (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur financier
    debut_mandat: 20/07/2007
    nom_de_famille: Lezeau
    nom: Michel Lezeau
    type: depute
  depute_267289:
    fonctions:
      - commission des affaires sociales / secrétaire / 
      - mission d'information commune sur l'indemnisation des victimes des maladies nosocomiales et accès au dossier médical / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 267289
    extras:
      - commission du fonds national pour l'archéologie préventive / membre titulaire
      - haut conseil des musées de france / membre suppléant
    adresses:
      - Hôtel de Ville 6 Rue Gambetta 45200 Montargis Téléphone : 02 38 95 10 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loiret (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Door
    place_hemicycle: 279
    autresmandats:
      - Maire de Montargis, Loiret (15022 habitants)
    mails:
      - doorjp@wanadoo.fr
      - jpdoor@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267289.asp
    profession: Cardiologue
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Door
    type: depute
  depute_267297:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des finances / secrétaire / 
    sexe: H
    id_an: 267297
    extras:
      - conseil d'administration de l'ecole nationale d'administration / membre titulaire
      - haut conseil du secteur public / membre titulaire
      - conseil d'administration de l'établissement public de réalisation de défaisance / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 62 91 Télécopie : 01 40 63 50 42 
      - Permanence 2 Rue Bayle de Seyches 47200 Marmande Téléphone : 05 53 89 31 85 Télécopie : 05 53 20 68 85 
    circonscription: Lot-et-Garonne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Diefenbacher
    place_hemicycle: 128
    mails:
      - mdiefenbacher@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267297.asp
    profession: Conseiller Maître à la Cour des comptes
    site_web: http://www.mdiefenbacher.org
    debut_mandat: 20/06/2007
    nom: Michel Diefenbacher
    type: depute
  depute_267306:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267306
    adresses:
      - 4 Place Jean-Antoine Pourtier 63890 Saint-Amant-Roche-Savine Téléphone : 04 73 95 74 90 Télécopie : 04 73 95 71 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Puy-de-Dôme (5ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Chassaigne
    place_hemicycle: 594
    autresmandats:
      - Maire de Saint-Amant-Roche-Savine, Puy-de-Dôme (531 habitants)
    mails:
      - chassaigne.a@wanadoo.fr
      - achassaigne@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267306.asp
    profession: Principal de collège
    site_web: http://www.andrechassaigne.org
    debut_mandat: 20/06/2007
    nom: André Chassaigne
    type: depute
  depute_267309:
    place_hemicycle: 370
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du conseil régional (Franche-Comté)
    sexe: H
    id_an: 267309
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267309.asp
    circonscription: Haute-Saône (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin
    debut_mandat: 19/04/2008
    nom_de_famille: Debray
    nom: Patrice Debray
    type: depute
  depute_267314:
    fonctions:
      - commission des finances / membre / 
    sexe: F
    id_an: 267314
    extras:
      - comité consultatif du secteur financier / membre titulaire
      - comité d'enquête sur le coût et le rendement des services publics / membre suppléante
    adresses:
      - Permanence parlementaire 110 Rue Aristide Briand BP 90112 72500 Château-du-Loir Téléphone : 02 43 44 46 97 Télécopie : 02 43 46 16 55 
      - Permanence parlementaire 11 Place Thiers 72200 La Flèche Téléphone : 02 43 94 75 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Sarthe (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Pavy
    place_hemicycle: 219
    autresmandats:
      - Vice-présidente de la communauté de communes Loir et Bercé
      - Maire de Saint-Pierre-de-Chevillé, Sarthe (342 habitants)
      - Membre du conseil général (Sarthe)
    mails:
      - bpavy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267314.asp
    profession: Comptable
    site_web: http://www.beatricepavy.blogspot.com
    debut_mandat: 20/06/2007
    nom: Béatrice Pavy
    type: depute
  depute_267317:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267317
    extras:
      - conseil d'administration de l'établissement public de sécurité ferroviaire / membre titulaire
    adresses:
      - 119 Rue de Malpalu "Résidence des Noisetiers" 72000 Le Mans Téléphone : 02 43 76 07 41 Télécopie : 02 43 76 12 79 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Sarthe (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Mèner
    place_hemicycle: 205
    autresmandats:
      - Membre du conseil général (Sarthe)
    mails:
      - dominique.le-mener@voila.fr
      - dlemener@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267317.asp
    profession: Juriste
    debut_mandat: 20/06/2007
    nom: Dominique Le Mèner
    type: depute
  depute_267324:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267324
    extras:
      - conseil d'administration de l'institut des hautes études pour la science et la technologie / membre titulaire
    adresses:
      - 5 Rue du Colonel Renard 88300 Neufchâteau Téléphone : 03 29 94 20 86 Télécopie : 03 29 94 35 13 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vosges (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gaultier
    place_hemicycle: 117
    autresmandats:
      - Vice-président du conseil général (Vosges)
    mails:
      - jjgaultier.depute@wanadoo.fr
      - jjgaultier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267324.asp
    profession: Médecin biologiste
    debut_mandat: 20/06/2007
    nom: Jean-Jacques Gaultier
    type: depute
  depute_267327:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267327
    adresses:
      - 4 Rue Georges Clemenceau 90000 Belfort Téléphone : 03 84 22 19 07 Télécopie : 03 84 28 36 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Territoire-de-Belfort (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Meslot
    place_hemicycle: 217
    autresmandats:
      - Membre du conseil général (Territoire de Belfort)
    mails:
      - dmeslot@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267327.asp
    profession: Cadre bancaire
    site_web: http://www.damienmeslot.com
    debut_mandat: 20/06/2007
    nom: Damien Meslot
    type: depute
  depute_267330:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 267330
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 9 Faubourg de Lyon 90000 Belfort Téléphone : 03 84 90 15 10 Télécopie : 03 84 90 15 35 
    circonscription: Territoire-de-Belfort (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Zumkeller
    place_hemicycle: 214
    autresmandats:
      - Maire de Valdoie, Territoire-de-Belfort (4843 habitants)
    mails:
      - michel.zumkeller@wanadoo.fr
      - mzumkeller@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267330.asp
    profession: Comptable
    site_web: http://www.michelzumkeller.net
    debut_mandat: 20/06/2007
    nom: Michel Zumkeller
    type: depute
  depute_267336:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267336
    adresses:
      - 10  Avenue de Vallouise 05120 L'Argentière-la-Bessée Téléphone : 04 92 21 33 81 Télécopie : 04 92 21 43 73 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hautes-Alpes (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Giraud
    place_hemicycle: 620
    autresmandats:
      - Vice-président du conseil régional (Provence-Alpes-Côte-d'Azur)
      - Maire de L'Argentière-la-Bessée, Hautes-Alpes (2289 habitants)
    mails:
      - jgiraud@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267336.asp
    profession: Administrateur civil hors-classe
    site_web: http://www.joelgiraud.net
    debut_mandat: 20/06/2007
    nom: Joël Giraud
    type: depute
  depute_267350:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 267350
    extras:
      - conseil national du tourisme / membre titulaire
    adresses:
      - 103 Boulevard Cassagnes 66140 Canet-en-Roussillon Téléphone : 04 68 80 25 63 Télécopie : 04 68 80 33 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie Place de l'Hôtel de Ville 66140 Canet-en-Roussillon 
    circonscription: Pyrénées-Orientales (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Franco
    place_hemicycle: 145
    autresmandats:
      - Maire de Canet-en-Roussillon, Pyrénées-Orientales (10182 habitants)
      - Vice-présidente de la communauté d'agglomération Têt Méditerranée
    mails:
      - arlette.franco@free.fr
      - afranco@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267350.asp
    profession: Enseignante
    debut_mandat: 20/06/2007
    nom: Arlette Franco
    type: depute
  depute_267355:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267355
    adresses:
      - Permanence 2 Rue du Docteur Bronner 67600 Sélestat Téléphone : 03 88 92 32 45 Télécopie : 03 88 82 84 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Herth
    place_hemicycle: 163
    autresmandats:
      - Membre du Conseil municipal d'Artolsheim, Bas-Rhin (723 habitants)
    mails:
      - aherth@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267355.asp
    profession: Agriculteur
    site_web: http://www.antoine-herth.fr
    debut_mandat: 20/06/2007
    nom: Antoine Herth
    type: depute
  depute_267358:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 267358
    extras:
      - conseil d'orientation de l'observatoire national sur les effets du réchauffement climatique en france métropolitaine et dans les départements et territoires d'outre-mer / membre titulaire
    adresses:
      - Mairie Place de l'Hôtel de Ville 68150 Ribeauvillé Téléphone : 03 89 73 20 00 Télécopie : 03 89 73 37 18 
      - Permanence parlementaire 10  Grand'Rue 68230 Turckheim Téléphone : 03 89 27 29 64 Télécopie : 03 89 27 16 73 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Christ
    place_hemicycle: 19
    autresmandats:
      - Maire de Ribeauvillé, Haut-Rhin (4929 habitants)
    mails:
      - christjl@wanadoo.fr
      - jlchrist@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267358.asp
    profession: Chef d'entreprise
    site_web: http://www.jlchrist-depute.com
    debut_mandat: 20/06/2007
    nom: Jean-Louis Christ
    type: depute
  depute_267378:
    fonctions:
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 267378
    extras:
      - comité national des retraités et des personnes âgées / membre titulaire
      - commission nationale consultative des droits de l'homme / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 52 Cours Lafayette 83000 Toulon Téléphone : 04 94 24 06 23 Télécopie : 04 94 24 91 01 
    circonscription: Var (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Levy
    place_hemicycle: 312
    autresmandats:
      - Première adjointe de Toulon, Var (160406 habitants)
    mails:
      - glevy@assemblee-nationale.fr
      - permanence.levy@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267378.asp
    profession: Expert foncier et commercial
    site_web: http://www.genevievelevy.com
    debut_mandat: 20/06/2007
    nom: Geneviève Levy
    type: depute
  depute_267382:
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267382
    extras:
      - commission nationale de la vidéosurveillance / membre titulaire
    adresses:
      - Mairie de Villemomble 13 Bis Rue d'Avron 93250 Villemomble Téléphone : 01 49 35 25 55 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Calméjane
    place_hemicycle: 31
    autresmandats:
      - Maire de Villemomble, Seine-Saint-Denis (26991 habitants)
    mails:
      - p.calmejane@mairie-villemomble.fr
      - pcalmejane@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267382.asp
    profession: Ingénieur
    debut_mandat: 20/06/2007
    nom: Patrice Calméjane
    type: depute
  depute_267399:
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 267399
    adresses:
      - 33 Rue Mignet 13100 Aix-en-Provence 
      - Mairie Place de l'Hôtel de Ville 13100 Aix-en-Provence Téléphone : 04 42 91 99 55 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (14ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Joissains-Masini
    place_hemicycle: 295
    autresmandats:
      - Maire d'Aix-en-Provence, Bouches-du-Rhône (134222 habitants)
    mails:
      - mjoissains@assemblee-nationale.fr
      - depute@marysejoissains.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267399.asp
    profession: Avocat
    site_web: http://www.marysejoissains.com
    debut_mandat: 20/06/2007
    nom: Maryse Joissains-Masini
    type: depute
  depute_267407:
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - assemblée nationale / secrétaire / 27/06/2007
      - commission des affaires étrangères / membre / 
      - délégation chargée de la communication audiovisuelle et de la presse / membre / 
      - délégation chargée de la communication et de la presse / membre / 
    sexe: H
    id_an: 267407
    adresses:
      - Hôtel du Département Rond-Point du Maréchal Leclerc 20405 Bastia cedex Téléphone : 04 95 55 55 51 Télécopie : 04 95 55 02 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Corse (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Giacobbi
    place_hemicycle: 616
    autresmandats:
      - Président du conseil général (Haute-Corse)
    mails:
      - pgiacobbi@cg2b.fr
      - pgiacobbi@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267407.asp
    profession: Administrateur civil hors classe au ministère de l'équipement
    site_web: http://www.paul-giacobbi.org
    debut_mandat: 20/06/2007
    nom: Paul Giacobbi
    type: depute
  depute_267424:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 267424
    extras:
      - commission de suivi de la détention provisoire / membre titulaire
    adresses:
      - Permanence parlementaire 3 Rue de la fontaine 33500 Pomerol Téléphone : 05 57 51 14 72 Télécopie : 05 57 51 77 41 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Garraud
    place_hemicycle: 6
    mails:
      - jpgarraud@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267424.asp
    profession: Magistrat
    site_web: http://www.jpgarraud.net
    debut_mandat: 20/06/2007
    nom: Jean-Paul Garraud
    type: depute
  depute_267429:
    place_hemicycle: 196
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 267429
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267429.asp
    mails:
      - dcinieri@assemblee-nationale.fr
    adresses:
      - Permanence 1 Rue Courbon-Brioude 42700 Firminy Téléphone : 04 77 89 20 44 Télécopie : 04 77 10 93 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.dinocinieri.com
    profession: Consultant sécurité
    debut_mandat: 20/06/2007
    nom_de_famille: Cinieri
    nom: Dino Cinieri
    type: depute
  depute_267433:
    place_hemicycle: 306
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Cholet, Maine-et-Loire (54198 habitants)
    sexe: H
    id_an: 267433
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267433.asp
    mails:
      - gbourdouleix@assemblee-nationale.fr
      - gbourdouleix@ville-cholet.fr
    adresses:
      - Permanence parlementaire 7  Rue Travot 49300 Cholet Téléphone : 02 41 70 03 51 Télécopie : 02 41 49 13 52 
      - Mairie Place Jean Moulin 49300 Cholet Téléphone : 02 41 49 25 08 Télécopie : 02 41 49 26 26 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 02 10 Télécopie : 01 40 63 02 90 
    circonscription: Maine-et-Loire (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chargé d'enseignement
    debut_mandat: 20/06/2007
    nom_de_famille: Bourdouleix
    nom: Gilles Bourdouleix
    type: depute
  depute_267440:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - commission des lois / membre / 
    sexe: H
    id_an: 267440
    extras:
      - comité consultatif des subventions aux exploitants d'aérodromes / membre titulaire
    adresses:
      - Permanence 7 Place de la République 13700 Marignane Téléphone : 04 42 77 14 73 Télécopie : 04 42 09 99 37 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 59 
      - Mairie Place des Droits de l'Homme 13960 Sausset-les-Pins Téléphone : 04 42 44 51 51 Télécopie : 04 42 44 62 96 
    circonscription: Bouches-du-Rhône (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Diard
    place_hemicycle: 234
    autresmandats:
      - Membre de la communauté urbaine Marseille Provence Métropole
      - Maire de Sausset-les-Pins, Bouches-du-Rhône (7233 habitants)
    mails:
      - ediard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267440.asp
    profession: Consultant en gestion
    site_web: http://www.ericdiard.fr
    debut_mandat: 20/06/2007
    nom: Éric Diard
    type: depute
  depute_267450:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / membre / 
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 267450
    adresses:
      - Permanence 81 Avenue Maréchal Lyautey 21000 Dijon 
    circonscription: Côte-d'Or (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Delatte
    place_hemicycle: 221
    autresmandats:
      - Maire de Saint-Apollinaire, Côte-d'Or (5016 habitants)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267450.asp
    mails:
      - permanence@remi-delatte.com
    site_web: http://www.remi-delatte.com
    profession: Agriculteur-propriétaire exploitant
    debut_mandat: 20/06/2007
    nom: Rémi Delatte
    type: depute
  depute_267457:
    place_hemicycle: 134
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Adjoint au Maire de Béziers, Hérault (69294 habitants)
    sexe: H
    id_an: 267457
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267457.asp
    circonscription: Hérault (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin cardiologue (Chef de service)
    debut_mandat: 04/07/2007
    nom_de_famille: Aboud
    nom: Élie Aboud
    type: depute
  depute_267459:
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - assemblée nationale / secrétaire / 27/06/2007
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléante / 
      - délégation chargée de l'application du statut du député / membre / 
      - commission des affaires culturelles et de l'éducation / secrétaire / 
      - délégation chargée de la communication audiovisuelle et de la presse / membre / 
      - délégation chargée de la communication et de la presse / membre / 
    sexe: F
    id_an: 267459
    extras:
      - conseil national du syndrome immunodéficitaire acquis / membre titulaire
      - conseil supérieur de la mutualité / membre titulaire
    adresses:
      - Permanence parlementaire 11 Place Saint-Denis 37400 Amboise Téléphone : 02 47 57 68 57 Télécopie : 02 47 57 74 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Indre-et-Loire (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Greff
    place_hemicycle: 263
    autresmandats:
      - Membre du conseil régional (Centre)
    mails:
      - c.greff@wanadoo.fr
      - cgreff@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267459.asp
    profession: Infirmière
    site_web: http://www.claudegreff.fr
    debut_mandat: 20/06/2007
    nom: Claude Greff
    type: depute
  depute_267469:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267469
    extras:
      - comité des finances locales / membre titulaire
    adresses:
      - Permanence, Place Saint-Pierre 3 Rue des Patenôtriers 49400 Saumur Téléphone : 02 41 67 65 26 Télécopie : 02 41 67 65 50 
      - Permanence, Mme Maryvonne Martin 2 Bis Rue J. du Bellay 49380 Thouarcé Téléphone : 02 41 78 34 33 Télécopie : 02 41 54 59 96 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Maine-et-Loire (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Piron
    place_hemicycle: 287
    autresmandats:
      - Membre du Conseil municipal de Thouarcé, Maine-et-Loire (1677 habitants)
      - Président de la communauté de communes des Coteaux-du-Layon
      - Membre du conseil général (Maine-et-Loire)
    mails:
      - michelpirondepute@wanadoo.fr
      - mpiron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267469.asp
    profession: Enseignant, puis chef d'entreprise
    site_web: http://www.michel-piron.fr
    debut_mandat: 20/06/2007
    nom: Michel Piron
    type: depute
  depute_267479:
    place_hemicycle: 473
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Maire de Saint-Pons-de-Thomières, Hérault (2287 habitants)
      - Président de la Communauté de communes du Pays Saint-Ponais
      - Membre du conseil général (Hérault)
    sexe: H
    id_an: 267479
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267479.asp
    mails:
      - kmesquida@assemblee-nationale.fr
      - mesquida.depute@wanadoo.fr
    adresses:
      - 1  Rue Général Thomières 34500 Béziers Téléphone : 04 67 11 29 61 Télécopie : 04 67 11 26 32 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hérault (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Ingénieur
    debut_mandat: 20/06/2007
    nom_de_famille: Mesquida
    nom: Kléber Mesquida
    type: depute
  depute_267492:
    fonctions:
      - commission de la défense nationale et des forces armées / secrétaire / 
    sexe: H
    id_an: 267492
    extras:
      - commission nationale pour l'élimination des mines antipersonnel / membre titulaire
    adresses:
      - Permanence Place Victor Brachelet 59490 Somain Téléphone : 03 27 98 82 21 Télécopie : 03 27 98 92 26 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (16ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Candelier
    place_hemicycle: 582
    autresmandats:
      - Président de la Communauté de communes de Coeur d'Ostrevent
      - Maire de Bruille-lez-Marchiennes, Nord (1213 habitants)
    mails:
      - jjcandelier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267492.asp
    profession: Retraité de la fonction publique
    site_web: http://www.jeanjacquescandelier.fr
    debut_mandat: 20/06/2007
    nom: Jean-Jacques Candelier
    type: depute
  depute_267499:
    fonctions:
      - commission de la défense nationale et des forces armées / secrétaire / 
    sexe: H
    id_an: 267499
    adresses:
      - Permanence parlementaire 108 Avenue Georges Clemenceau Bât.C3 69230 Saint-Genis-Laval Téléphone : 04 72 39 94 09 Télécopie : 04 72 39  96 51 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Guilloteau
    place_hemicycle: 349
    autresmandats:
      - Membre du conseil général (Rhône)
    mails:
      - cguilloteau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267499.asp
    profession: Ancien assistant parlementaire
    site_web: http://www.christopheguilloteau.com
    debut_mandat: 20/06/2007
    nom: Christophe Guilloteau
    type: depute
  depute_267506:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission de la défense nationale et des forces armées / vice-président / 
    sexe: H
    id_an: 267506
    extras:
      - comité de surveillance de la caisse d'amortissement de la dette sociale / membre titulaire
      - conseil d'administration de l'institut des hautes études de défense nationale / membre titulaire
    adresses:
      - Le Concorde 280 Avenue Maréchal Foch 83000 Toulon Téléphone : 04 94 24 42 19 Télécopie : 04 94 24 12 34 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Var (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Vitel
    place_hemicycle: 327
    autresmandats:
      - Vice-président du conseil général (Var)
    mails:
      - vitel.depute@wanadoo.fr
      - pvitel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267506.asp
    profession: Chirurgien plasticien
    site_web: http://www.philippevitel.com
    debut_mandat: 20/06/2007
    nom: Philippe Vitel
    type: depute
  depute_267512:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267512
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 8 Rue Lamartine 12400 Saint-Affrique Téléphone : 05 65 99 05 81 Télécopie : 05 65 49 38 65 
    circonscription: Aveyron (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Marc
    place_hemicycle: 30
    autresmandats:
      - Premier Vice-président du conseil général (Aveyron)
    mails:
      - amarc@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267512.asp
    profession: Retraité de l'enseignement
    site_web: http://www.alainmarc.com
    debut_mandat: 20/06/2007
    nom: Alain Marc
    type: depute
  depute_267519:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267519
    extras:
      - observatoire national de la sécurité des établissements scolaires et d'enseignement supérieur / membre suppléant
    adresses:
      - Mairie 30000 Nîmes Téléphone : 04 66 76 51 05 Télécopie : 04 66 76 51 36 
      - 35 Avenue Georges Pompidou 30000 Nîmes Téléphone : 04 66 02 11 50 Télécopie : 04 66 02 43 32 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gard (1ère)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Lachaud
    place_hemicycle: 384
    autresmandats:
      - Adjoint au Maire de Nîmes, Gard (133424 habitants)
      - Vice-président de la communauté d'agglomération de Nîmes Métropole
    mails:
      - ylachaud@assemblee-nationale.fr
      - info@yvan-lachaud.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267519.asp
    profession: Chef d'établissement scolaire
    site_web: http://www.yvan-lachaud.com.
    debut_mandat: 20/06/2007
    nom: Yvan Lachaud
    type: depute
  depute_267527:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267527
    extras:
      - conseil national pour le développement, l'aménagement et la protection de la montagne / membre titulaire
      - conseil national des transports / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 111  Rue du Pont Immeuble "La Résidence" 74130 Bonneville Téléphone : 04 50 25 24 13 Télécopie : 04 50 25 95 83 
    circonscription: Haute-Savoie (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Saddier
    place_hemicycle: 231
    autresmandats:
      - Maire de Bonneville, Haute-Savoie (13000 habitants)
    mails:
      - msaddier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267527.asp
    profession: Cadre à la Chambre d'agriculture d'Annecy
    site_web: http://www.martial-saddier.fr
    debut_mandat: 20/06/2007
    nom: Martial Saddier
    type: depute
  depute_267532:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 267532
    adresses:
      - BP 64 74502 Évian-les-Bains cedex Téléphone : 04 50 83 10 07 Télécopie : 04 50 75 68 85 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 02 63 Télécopie : 01 40 63 02 93 
      - Représentation parlementaire 5 Rue de l'Hôtel de Ville 74200 Thonon-les-Bains Téléphone : 04 50 70 12 19 Télécopie : 04 50 71 70 19 
    circonscription: Haute-Savoie (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Francina
    place_hemicycle: 126
    autresmandats:
      - Maire d'Évian-les-Bains, Haute-Savoie (7273 habitants)
    mails:
      - mfrancina@assemblee-nationale.fr
      - p.mahut@marcfrancina.net
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267532.asp
    profession: Conseiller financier et bancaire
    site_web: http://www.marcfrancina.net
    debut_mandat: 20/06/2007
    nom: Marc Francina
    type: depute
  depute_267542:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 267542
    extras:
      - conseil supérieur de l'établissement national des invalides de la marine / membre titulaire
    adresses:
      - 1 Rue des Carmélites 22200 Guingamp Téléphone : 02 96 40 08 97 Télécopie : 02 96 44 26 09 
      - Hôtel de Ville 1 Place de la Mairie 22340 Treffrin 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côtes-d'Armor (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Oget
    place_hemicycle: 436
    autresmandats:
      - Maire de Treffrin, Côtes-d'Armor (572 habitants)
    mails:
      - mroget@assemblee-nationale.fr
      - oget.mr@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267542.asp
    profession: Directrice d'association
    debut_mandat: 20/06/2007
    nom: Marie-Renée Oget
    type: depute
  depute_267545:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / secrétaire / 
    sexe: F
    id_an: 267545
    adresses:
      - Permanence parlementaire 27 B Rue Clément Marot 25000 Besançon Téléphone : 03 81 21 24 25 Télécopie : 03 81 83 49 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Doubs (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Branget
    place_hemicycle: 8
    autresmandats:
      - Membre du Conseil municipal de Besançon, Doubs (117696 habitants)
    mails:
      - francoise@branget.com
      - fbranget@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267545.asp
    profession: Gestionnaire en immobilier
    site_web: http://www.branget.com
    debut_mandat: 20/06/2007
    nom: Françoise Branget
    type: depute
  depute_267551:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 267551
    adresses:
      - 13 Place Leopold 54300 Lunéville Téléphone : 03 83 73 79 58 Télécopie : 03 83 73 78 02 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meurthe-et-Moselle (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lamblin
    place_hemicycle: 38
    autresmandats:
      - Maire de Lunéville, Meurthe-et-Moselle (20199 habitants)
    mails:
      - permanence.lamblin@yahoo.fr
      - jlamblin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267551.asp
    profession: Vétérinaire
    site_web: http://www.jacqueslamblin.fr
    debut_mandat: 20/06/2007
    nom: Jacques Lamblin
    type: depute
  depute_267556:
    place_hemicycle: 317
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Sarrebourg, Moselle (13341 habitants)
    sexe: H
    id_an: 267556
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267556.asp
    mails:
      - a.marty-depute@wanadoo.fr
      - amarty@assemblee-nationale.fr
    adresses:
      - 16 Rue de la Gare 57400 Sarrebourg Téléphone : 03 87 25 74 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville Avenue du Général de Gaulle 57400 Sarrebourg Téléphone : 03 87 03 05 06 Télécopie : 03 87 03 05 19 
    circonscription: Moselle (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Gynécologue obstétricien
    debut_mandat: 20/06/2007
    nom_de_famille: Marty
    nom: Alain Marty
    type: depute
  depute_267561:
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 267561
    adresses:
      - 4 Rue Armand Cambon 82000 Montauban Téléphone : 05 63 20 40 83 Télécopie : 05 63 63 96 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Tarn-et-Garonne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Barèges
    place_hemicycle: 188
    autresmandats:
      - Maire de Montauban, Tarn-et-Garonne (51855 habitants)
    mails:
      - brigitte.bareges@wanadoo.fr
      - bbareges@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267561.asp
    profession: Avocat
    site_web: http://www.brigittebareges.com
    debut_mandat: 20/06/2007
    nom: Brigitte Barèges
    type: depute
  depute_267570:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267570
    extras:
      - conseil de surveillance du fonds de financement de la protection complémentaire  de la couverture universelle du risque maladie / membre titulaire
    adresses:
      - Permanence 44 Rue du Général de Gaulle 89270 Vermenton Téléphone : 03 86 31 91 80 Télécopie : 03 86 31 91 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yonne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Rolland
    place_hemicycle: 300
    autresmandats:
      - Membre du Conseil municipal de Vermenton, Yonne (1199 habitants)
      - Président de la communauté de communes entre Cure et Yonne
      - Président du conseil général (Yonne)
    mails:
      - jeanmarie.rolland@free.fr
      - jmrolland@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267570.asp
    profession: Médecin généraliste
    debut_mandat: 20/06/2007
    nom: Jean-Marie Rolland
    type: depute
  depute_267573:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267573
    adresses:
      - Mairie 2 Rue Sérafini 20000 Ajaccio Téléphone : 04 95 21 18 92 Télécopie : 04 95 21 54 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 2 Rue du Docteur Versini 20000 Ajaccio Téléphone : 04 95 21 89 54 Télécopie : 04 95 22 16 93 
    circonscription: Corse-du-Sud (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Renucci
    place_hemicycle: 464
    autresmandats:
      - Maire d'Ajaccio, Corse-du-Sud (52880 habitants)
    mails:
      - srenucci@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267573.asp
    profession: Pédiatre
    site_web: http://simon-renucci.org
    debut_mandat: 20/06/2007
    nom: Simon Renucci
    type: depute
  depute_267576:
    place_hemicycle: 228
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission des lois / membre / 
    sexe: H
    id_an: 267576
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267576.asp
    mails:
      - marcelbonnot@yahoo.fr
      - mbonnot@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 1  Rue de la Schliffe BP 67361 25207 Montbéliard cedex Téléphone : 03 81 91 84 60 Télécopie : 03 81 91 79 95 
    circonscription: Doubs (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Bonnot
    nom: Marcel Bonnot
    type: depute
  depute_267585:
    fonctions:
      - commission des affaires européennes / secrétaire / 
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267585
    adresses:
      - Permanence parlementaire 69  Rue du Général Leclerc BP 70707 59510 Hem Téléphone : 03 20 45 48 48 Télécopie : 03 20 02 28 04 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie Rue du Général Leclerc 59510 Hem Téléphone : 03 20 66 58 00 Télécopie : 03 20 81 17 18 
    circonscription: Nord (7ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Vercamer
    place_hemicycle: 377
    autresmandats:
      - Maire de Hem, Nord (19675 habitants)
    mails:
      - fvercamer@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267585.asp
    profession: Ingénieur
    site_web: http://www.vercamer.fr
    debut_mandat: 20/06/2007
    nom: Francis Vercamer
    type: depute
  depute_267598:
    place_hemicycle: 314
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Vice-présidente du conseil général (Var)
    sexe: F
    id_an: 267598
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267598.asp
    circonscription: Var (6ème)
    adresses:
      - 13  Rue Victor Hugo 83270 Saint Cyr sur Mer Téléphone : 04 94 26 18 37 Télécopie : 04 94 26 17 40 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.josettepons.fr
    debut_mandat: 20/06/2007
    nom_de_famille: Pons
    nom: Josette Pons
    type: depute
  depute_267606:
    place_hemicycle: 392
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Membre du Conseil municipal de Lévis-Saint-Nom, Yvelines (1696 habitants)
      - Vice-président du conseil général (Yvelines)
    sexe: H
    id_an: 267606
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267606.asp
    circonscription: Yvelines (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Professeur agrégé de géographie
    debut_mandat: 20/07/2007
    nom_de_famille: Vandewalle
    nom: Yves Vandewalle
    type: depute
  depute_267622:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 267622
    extras:
      - commission nationale de la vidéosurveillance / membre titulaire
    adresses:
      - Permanence parlementaire 35 Rue de Paris 91100 Corbeil-Essonnes Téléphone : 01 60 88 01 23 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Essonne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Valls
    place_hemicycle: 425
    autresmandats:
      - Maire d'Évry, Essonne (48952 habitants)
    mails:
      - mvalls@assemblee-nationale.fr
      - maire@mairie-evry.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267622.asp
    profession: Conseiller en communication
    site_web: http://www.valls.fr
    debut_mandat: 20/06/2007
    nom: Manuel Valls
    type: depute
  depute_267641:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267641
    adresses:
      - Permanence 3 Rue rue Lamarque BP 30 18201 Saint-Amand-Montrond  Téléphone : 02 48 96 09 44 Télécopie : 02 48 60 18 95 
      - Mairie Place des Ormes 18130 Dun-sur-Auron Téléphone : 02 48 66 64 20 Télécopie : 02 48 59 84 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Cher (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cosyns
    place_hemicycle: 296
    autresmandats:
      - Maire de Dun-sur-Auron, Cher (4010 habitants)
      - Membre de la communauté de communes du Dunois
    mails:
      - lcosyns@assemblee-nationale.fr
      - l.cosyns.sam@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267641.asp
    profession: Agent général d'assurances
    site_web: http://www.louiscosyns.fr
    debut_mandat: 20/06/2007
    nom: Louis Cosyns
    type: depute
  depute_267644:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 267644
    extras:
      - commission nationale de concertation sur les risques miniers / membre titulaire
      - conseil d'orientation pour la prévention des risques naturels majeurs / membre titulaire
    adresses:
      - Permanence parlementaire 15 Bis Route de Dijon 21600 Longvic Téléphone : 03 80 65 87 87 Télécopie : 03 80 65 87 88 
      - Mairie 21600 Longvic Téléphone : 03 80 68 44 00 Télécopie : 03 80 68 44 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côte-d'Or (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Darciaux
    place_hemicycle: 460
    autresmandats:
      - Maire de Longvic, Côte-d'Or (8962 habitants)
      - Membre de la communauté de l'agglomération dijonnaise
    mails:
      - cadarciaux@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267644.asp
    profession: Enseignante
    debut_mandat: 20/06/2007
    nom: Claude Darciaux
    type: depute
  depute_267647:
    place_hemicycle: 15
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire du Grau-du-Roi, Gard (8000 habitants)
    sexe: H
    id_an: 267647
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267647.asp
    mails:
      - emourrut.depute@wanadoo.fr
      - emourrut@assemblee-nationale.fr
    adresses:
      - Permanence 22 Rue de la Poissonnerie BP 200 30240 Le Grau-du-Roi Téléphone : 04 66 51 73 64 Télécopie : 04 66 51 88 37 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gard (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Commerçant retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Mourrut
    nom: Étienne Mourrut
    type: depute
  depute_267650:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 267650
    extras:
      - conseil d'administration de la société nationale de programme radio france internationale (rfi) / membre titulaire
    adresses:
      - Hôtel de Ville 30400 Villeneuve-lèz-Avignon Téléphone : 04 90 27 49 04 Télécopie : 04 90 27 49 79 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gard (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Roubaud
    place_hemicycle: 302
    autresmandats:
      - Vice-président de la communauté d'agglomération du Grand Avignon (COGA)
      - Maire de Villeneuve-lès-Avignon, Gard (12500 habitants)
    mails:
      - jmroubaud@assemblee-nationale.fr
      - permanencejmroubaud@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267650.asp
    profession: Pharmacien
    site_web: http://www.jmroubaud.com
    debut_mandat: 20/06/2007
    nom: Jean-Marc Roubaud
    type: depute
  depute_267662:
    place_hemicycle: 356
    fonctions:
      - commission des affaires étrangères / secrétaire / 
    autresmandats:
      - Maire de Vienne, Isère (29972 habitants)
    sexe: H
    id_an: 267662
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267662.asp
    mails:
      - jremiller@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville, Cabinet du Maire 1 Place de l'Hôtel de Ville BP 126 38209 Vienne cedex Téléphone : 04 74 78 30 00 (Standard) Téléphone : 04 74 78 30 15 (Cabinet) Télécopie : 04 74 31 78 67 
      - Permanence parlementaire 21 Place Charles de Gaulle BP 134 38209 Vienne cedex Téléphone : 04 74 59 29 55 Télécopie : 04 74 78 22 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre bancaire retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Remiller
    nom: Jacques Remiller
    type: depute
  depute_267673:
    fonctions:
      - commission de la défense nationale et des forces armées / vice-président / 
    sexe: H
    id_an: 267673
    extras:
      - conseil supérieur de la réserve militaire / membre suppléant
    adresses:
      - Permanence 3  Boulevard des Lices 81100 Castres Téléphone : 05 63 71 29 23 Télécopie : 05 63 59 82 71 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Tarn (3ème)
    groupe:
      - nouveau centre / apparenté
    nom_de_famille: Folliot
    place_hemicycle: 387
    autresmandats:
      - Membre du Conseil municipal de Castres, Tarn (43454 habitants)
    mails:
      - pfolliot@assemblee-nationale.fr
      - contact@philippe-folliot.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267673.asp
    profession: Directeur d'un organisme de financement du logement social
    site_web: http://www.philippe-folliot.fr
    debut_mandat: 20/06/2007
    nom: Philippe Folliot
    type: depute
  depute_267689:
    place_hemicycle: 33
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Président de l'Assemblée de Corse
    sexe: H
    id_an: 267689
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267689.asp
    mails:
      - cderoccaserra@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 2 Rue Joseph Pietri 20137 Porto-Vecchio Téléphone : 04 95 23 30 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Corse-du-Sud (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.camillederoccaserra.com
    debut_mandat: 20/06/2007
    nom_de_famille: Serra
    nom: Camille de Rocca Serra
    type: depute
  depute_267695:
    fonctions:
      - commission de la défense nationale et des forces armées / vice-présidente / 
    sexe: F
    id_an: 267695
    extras:
      - conseil supérieur de la réserve militaire / membre titulaire
    adresses:
      - Permanence 43 D Rue Branda BP 21041 29210 Brest cedex 1 Téléphone : 02 98 33 21 80 Télécopie : 02 98 33 21 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Finistère (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Adam
    place_hemicycle: 424
    autresmandats:
      - Membre du conseil général (Finistère)
    mails:
      - patricia.adam-deputee@wanadoo.fr
      - padam@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267695.asp
    profession: Cadre d'action sociale
    debut_mandat: 20/06/2007
    nom: Patricia Adam
    type: depute
  depute_267698:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: F
    id_an: 267698
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
    adresses:
      - Téléphone mobile : 06 63 34 34 97 Téléphone mobile : 06 61 32 10 48  marguerite.lamour@wanadoo.fr
      - Mairie Place André Colin 29830 Ploudalmézeau Téléphone : 02 98 48 02 56 Télécopie : 02 98 38 13 17 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 76 02 Télécopie : 01 40 63 78 43 
      - 6 Rue de Kerjolys 29830 Ploudalmézeau Téléphone : 02 98 48 14 99 Télécopie : 02 98 38 13 73 
    circonscription: Finistère (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lamour
    place_hemicycle: 129
    autresmandats:
      - Vice-présidente de la communauté de communes du Pays d'Iroise
      - Maire de Ploudalmézeau, Finistère (6087 habitants)
    mails:
      - mlamour@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267698.asp
    profession: Assistante administrative
    debut_mandat: 20/06/2007
    nom: Marguerite Lamour
    type: depute
  depute_267705:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission du développement durable et de l'aménagement du territoire / vice-président / 
    sexe: H
    id_an: 267705
    extras:
      - conseil d'orientation de l'observatoire national sur les effets du réchauffement climatique en france métropolitaine et dans les départements et territoires d'outre-mer / membre suppléant
    adresses:
      - Permanence 29 D Avenue du Bois Labbé 35000 Rennes Téléphone : 02 99 55 80 84 Télécopie : 02 99 55 18 28 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 74 57 
    circonscription: Ille-et-Vilaine (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Tourtelier
    place_hemicycle: 552
    mails:
      - ptourtelier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267705.asp
    profession: Professeur retraité
    site_web: http://www.philippe-tourtelier.fr
    debut_mandat: 20/06/2007
    nom: Philippe Tourtelier
    type: depute
  depute_267711:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 267711
    extras:
      - conseil national de l'enseignement supérieur et de la recherche / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 83  Rue Saint-Georges 54000 Nancy Téléphone : 03 83 35 57 21 Télécopie : 03 83 35 07 13 
    circonscription: Meurthe-et-Moselle (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Hénart
    place_hemicycle: 345
    autresmandats:
      - Adjoint au Maire de Nancy, Meurthe-et-Moselle (103606 habitants)
      - Membre de la communauté urbaine du Grand Nancy
    mails:
      - lhenart@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267711.asp
    profession: Juriste d'entreprise
    site_web: http://www.laurenthenart.com
    debut_mandat: 20/06/2007
    nom: Laurent Hénart
    type: depute
  depute_267719:
    place_hemicycle: 76
    fonctions:
      - délégation chargée d'examiner la recevabilité des propositions de loi / questeur, membre / 
      - commission des affaires sociales / membre / 
      - assemblée nationale / questeur / 27/06/2007
      - délégation chargée des activités internationales / questeur, membre / 
    sexe: H
    id_an: 267719
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267719.asp
    mails:
      - mallie.richard@wanadoo.fr
      - rmallie@assemblee-nationale.fr
    adresses:
      - 20 Rue Jules Ferry 13120 Gardanne Téléphone : 04 42 65 44 44 Télécopie : 04 42 65 44 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.depute-mallie.com
    profession: Docteur en chirurgie dentaire
    debut_mandat: 20/06/2007
    nom_de_famille: Mallié
    nom: Richard Mallié
    type: depute
  depute_267728:
    place_hemicycle: 304
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 267728
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre suppléant
      - conseil supérieur de l'énergie / membre suppléant
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267728.asp
    mails:
      - christophepriou@wanadoo.fr
      - cpriou@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 3  Rue du Beausoleil 44350 Guérande Téléphone : 02 40 62 02 72 Télécopie : 02 40 62 00 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre de chambre de commerce et d'industrie 
    debut_mandat: 20/06/2007
    nom_de_famille: Priou
    nom: Christophe Priou
    type: depute
  depute_267743:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267743
    extras:
      - commission nationale pour l'autonomie des jeunes / membre titulaire
    adresses:
      - 45   Rue du Pont de Pierre 60600 Clermont Téléphone : 03 44 19 07 87 Télécopie : 03 44 19 07 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Courtial
    place_hemicycle: 41
    autresmandats:
      - Maire d'Agnetz, Oise (2637 habitants)
    mails:
      - contact@edouard-courtial.org
      - ecourtial@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267743.asp
    profession: Consultant
    site_web: http://www.edouardcourtial.fr
    debut_mandat: 20/06/2007
    nom: Édouard Courtial
    type: depute
  depute_267762:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267762
    adresses:
      - Permanence 11 Place du Marché-aux-Fruits 59630 Bourbourg Téléphone : 03 28 22 33 33 Télécopie : 03 28 20 00 86 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie 59630 Brouckerque Téléphone : 03 28 27 12 00 Télécopie : 03 28 27 16 14 
    circonscription: Nord (14ème)
    groupe:
      - union pour un mouvement populaire / apparenté
    nom_de_famille: Decool
    place_hemicycle: 35
    autresmandats:
      - Membre du conseil général (Nord)
      - Maire de Brouckerque, Nord (1165 habitants)
    mails:
      - jpdecool@assemblee-nationale.fr
      - jpdecool@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267762.asp
    profession: Professeur
    site_web: http://www.jeanpierredecool.com
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Decool
    type: depute
  depute_267765:
    place_hemicycle: 67
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Premier vice-président de la communauté d'agglomération de Cambrai
      - Maire de Cambrai, Nord (33738 habitants)
    sexe: H
    id_an: 267765
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267765.asp
    mails:
      - fxvillain@assemblee-nationale.fr
      - fxvillain@wanadoo.fr
    adresses:
      - Hôtel de Ville 2 Rue de Nice 59400 Cambrai Téléphone : 03 27 73 21 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (18ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Villain
    nom: François-Xavier Villain
    type: depute
  depute_267768:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267768
    adresses:
      - 7  Rue du Maréchal Leclerc 59220 Denain Téléphone : 03 27 22 93 84 Télécopie : 03 27 22 93 87 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (19ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Roy
    place_hemicycle: 550
    autresmandats:
      - Maire de Denain, Nord (20356 habitants)
    mails:
      - proy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267768.asp
    profession: Enseignant
    site_web: http://www.patrick-roy.fr
    debut_mandat: 20/06/2007
    nom: Patrick Roy
    type: depute
  depute_267773:
    place_hemicycle: 5
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Membre du conseil général (Oise)
    sexe: H
    id_an: 267773
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267773.asp
    circonscription: Oise (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Agriculteur
    debut_mandat: 20/07/2007
    nom_de_famille: Patria
    nom: Christian Patria
    type: depute
  depute_267775:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 267775
    adresses:
      - Permanence 3 Place Charles de Gaulle 69130 Ecully 
      - Permanence 13 Rue Jean Moulin BP 101 69300 Caluire-et-Cuire Téléphone : 04 72 27 17 56 Télécopie : 04 78 08 51 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cochet
    place_hemicycle: 271
    autresmandats:
      - Maire de Caluire-et-Cuire, Rhône (41233 habitants)
    mails:
      - pcochet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267775.asp
    profession: Gérant de société
    site_web: http://www.philippecochet.com
    debut_mandat: 20/06/2007
    nom: Philippe Cochet
    type: depute
  depute_267787:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 267787
    extras:
      - conseil d'administration de la société nationale de programme réseau france-outre-mer (rfo) / membre titulaire
    adresses:
      - 14 Rue de la victoire 97400 Saint-Denis Téléphone : 02 62 30 60 60 Télécopie : 02 62 30 60 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Réunion (1ère)
    groupe:
      - union pour un mouvement populaire / apparenté
    nom_de_famille: Victoria
    place_hemicycle: 307
    autresmandats:
      - Membre du Conseil municipal de Saint-Denis, Réunion (132338 habitants)
    mails:
      - rpvictoria@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267787.asp
    profession: Directeur d'école
    site_web: http://www.rpvictoria.fr
    debut_mandat: 20/06/2007
    nom: René-Paul Victoria
    type: depute
  depute_267794:
    fonctions:
      - commission des affaires culturelles et de l'éducation / présidente / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: F
    id_an: 267794
    extras:
      - comité de suivi de l'agence française de l'adoption / membre titulaire
      - haut conseil de la famille / membre titulaire
      - conseil supérieur de l'adoption / membre titulaire
      - conseil supérieur de l' administration pénitentiaire / membre titulaire
    adresses:
      - Mairie 20 Boulevard Sadi Carnot 06110 Le Cannet Téléphone : 04 92 18 21 00 Télécopie : 04 92 18 21 01 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Alpes-Maritimes (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Tabarot
    place_hemicycle: 98
    autresmandats:
      - Maire du Cannet, Alpes-Maritimes (41885 habitants)
    mails:
      - mtabarot@assemblee-nationale.fr
      - 9circonscription@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267794.asp
    profession: Chef d'entreprise
    site_web: http://www.michele-tabarot.fr
    debut_mandat: 20/06/2007
    nom: Michèle Tabarot
    type: depute
  depute_267797:
    fonctions:
      - commission des affaires économiques / membre / 
      - délégation chargée de la communication et de la presse / présidente / 
      - assemblée nationale / vice-présidente / 26/09/2008
    sexe: F
    id_an: 267797
    extras:
      - conseil de surveillance du fonds de financement de l'allocation personnalisée d'autonomie / membre titulaire
    adresses:
      - Permanence 8 Rue de Venise 51100 Reims Téléphone : 03 26 82 42 15 Télécopie : 03 26 35 89 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Marne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Vautrin
    place_hemicycle: 82
    autresmandats:
      - Membre du Conseil municipal de Reims, Marne (187201 habitants)
    mails:
      - contact@catherine-vautrin.fr
      - cvautrin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267797.asp
    profession: Directeur marketing
    site_web: http://www.catherine-vautrin.fr
    debut_mandat: 20/06/2007
    nom: Catherine Vautrin
    type: depute
  depute_267810:
    place_hemicycle: 104
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Membre du conseil régional (Ile-de-France)
    sexe: F
    id_an: 267810
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267810.asp
    mails:
      - cbrunel@assemblee-nationale.fr
    adresses:
      - 6 Rue Konrad Adenauer  77600 Bussy Saint-Georges Téléphone : 01 60 06 35 27 Télécopie : 01 60 06 58 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-et-Marne (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.chantalbrunel.fr
    debut_mandat: 20/06/2007
    nom_de_famille: Brunel
    nom: Chantal Brunel
    type: depute
  depute_267813:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des lois / vice-président / 
    sexe: H
    id_an: 267813
    extras:
      - conseil d'administration de l'agence de l'environnement et de la maîtrise de l'énergie / membre titulaire
      - comité des finances locales / membre suppléant
      - conseil d'administration de l'institut national des hautes études de sécurité / membre titulaire
      - commission de surveillance et de contrôle des publications destinées à l'enfance et à l'adolescence / membre titulaire
    adresses:
      - Mairie de Combs-La-Ville Place de l'Hôtel de Ville 77385 Combs-la-Ville Cedex Téléphone : 01 64 13 16 03 Télécopie : 01 64 88 61 66 
      - 2  Avenue Victor Hugo 77170 Brie-Comte-Robert Téléphone : 01 60 62 24 21 Télécopie : 01 60 34 99 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-et-Marne (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Geoffroy
    place_hemicycle: 198
    autresmandats:
      - Maire de Combs-la-Ville, Seine-et-Marne (20953 habitants)
    mails:
      - geoffroy.depute@wanadoo.fr
      - ggeoffroy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267813.asp
    profession: Proviseur
    site_web: http://www.guy-geoffroy.com
    debut_mandat: 20/06/2007
    nom: Guy Geoffroy
    type: depute
  depute_267822:
    fonctions:
      - commission des lois / vice-président / 
    sexe: H
    id_an: 267822
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 29 Rue du Général de Gaulle 94430 Chennevières-sur-Marne Téléphone : 01 49 82 02 21 
    circonscription: Val-de-Marne (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bénisti
    place_hemicycle: 288
    autresmandats:
      - Maire de Villiers-sur-Marne, Val-de-Marne (26532 habitants)
    mails:
      - jabenisti@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267822.asp
    profession: Cadre d'entreprise
    site_web: http://www.jabenisti.com
    debut_mandat: 20/06/2007
    nom: Jacques Alain Bénisti
    type: depute
  depute_267827:
    place_hemicycle: 86
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Membre du Conseil municipal de Nogent-sur-Marne, Val-de-Marne (28191 habitants)
    sexe: F
    id_an: 267827
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267827.asp
    mails:
      - mamontchamp@assemblee-nationale.fr
    adresses:
      - Permanence 4 Rue Pasteur 94130 Nogent-sur-Marne Téléphone : 01 43 94 14 14 Télécopie : 01 40 63 63 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.marie-anne-montchamp.fr
    debut_mandat: 20/06/2007
    nom_de_famille: Montchamp
    nom: Marie-Anne Montchamp
    type: depute
  depute_267835:
    fonctions:
      - commission des affaires économiques / membre / 
      - mission d'information commune sur l'évaluation des dispositifs fiscaux d'encouragement à l'investissement locatif / membre / 
    sexe: H
    id_an: 267835
    extras:
      - conseil national de l'habitat / membre suppléant
      - commission nationale chargée de l'examen du respect des obligations de réalisation de logements sociaux / membre titulaire
      - conseil d'orientation de l'observatoire national des zones urbaines sensibles / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (11ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bouillonnec
    place_hemicycle: 452
    autresmandats:
      - Vice-président de la communauté d'agglomération du Val de Bièvre
      - Maire de Cachan, Val-de-Marne (24886 habitants)
    mails:
      - jylebouillonnec@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267835.asp
    profession: Avocat
    site_web: http://www.le-bouillonnec.net
    debut_mandat: 20/06/2007
    nom: Jean-Yves Le Bouillonnec
    type: depute
  depute_267859:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267859
    extras:
      - conseil de surveillance du fonds de financement de la protection complémentaire  de la couverture universelle du risque maladie / membre titulaire
    adresses:
      - Permanence parlementaire 39 Boulevard Rabelais 34000 Montpellier Téléphone : 04 67 54 33 94 Télécopie : 04 67 60 38 28 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hérault (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Domergue
    place_hemicycle: 130
    autresmandats:
      - Membre du conseil régional (Languedoc-Roussillon)
    mails:
      - jdomergue@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267859.asp
    profession: Chirurgien
    site_web: http://www.jacquesdomergue.com
    debut_mandat: 20/06/2007
    nom: Jacques Domergue
    type: depute
  depute_267862:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 267862
    adresses:
      - Permanence parlementaire 1  Boulevard du général Leclerc 34700 Lodève Téléphone : 04 67 88 61 21 Télécopie : 04 67 44 33 05 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hérault (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Lecou
    place_hemicycle: 212
    autresmandats:
      - Membre du Conseil municipal de Lodève, Hérault (6900 habitants)
    mails:
      - rlecou@assemblee-nationale.fr
      - permanence.lecou@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267862.asp
    profession: Cadre territorial
    site_web: http://www.robert-lecou.fr
    debut_mandat: 20/06/2007
    nom: Robert Lecou
    type: depute
  depute_267875:
    place_hemicycle: 303
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Président de la communauté d'agglomération des Hauts de Bièvre
      - Maire de Châtenay-Malabry, Hauts-de-Seine (32310 habitants)
    sexe: H
    id_an: 267875
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267875.asp
    circonscription: Hauts-de-Seine (13ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur de société
    debut_mandat: 05/01/2009
    nom_de_famille: Siffredi
    nom: Georges Siffredi
    type: depute
  depute_267886:
    fonctions:
      - commission des affaires étrangères / président / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: H
    id_an: 267886
    adresses:
      - Permanence parlementaire BP 80002 Cergy 95001 Cergy-Pontoise Cedex Téléphone : 01 34 69 17 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Poniatowski
    place_hemicycle: 285
    autresmandats:
      - Président de la communauté de communes de la Vallée de l'Oise et des Trois-Forêts
      - Maire de L'Isle-Adam, Val-d'Oise (11173 habitants)
    mails:
      - aponiatowski@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267886.asp
    profession: Directeur de société
    site_web: http://www.axelponiatowski.com
    debut_mandat: 20/06/2007
    nom: Axel Poniatowski
    type: depute
  depute_267895:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 267895
    extras:
      - conseil d'orientation de la simplification administrative / membre suppléant
    adresses:
      - 47 Rue de la Mairie 95330 Domont Téléphone : 01 39 35 55 01 Télécopie : 01 39 91 32 77 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Chartier
    place_hemicycle: 95
    autresmandats:
      - Maire de Domont, Val-d'Oise (14882 habitants)
    mails:
      - jchartier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267895.asp
    profession: Ancien associé gérant
    site_web: http://www.jeromechartier.fr
    debut_mandat: 20/06/2007
    nom: Jérôme Chartier
    type: depute
  depute_267903:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 267903
    extras:
      - comité de suivi de la mise en oeuvre des dispositions relatives au cinéma et autres arts et industries de l'image animée / membre suppléante
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 18 Boulevard Joseph Garnier 06000 Nice Téléphone : 04 93 52 34 80 Télécopie : 04 93 52 19 80 
    circonscription: Alpes-Maritimes (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Marland-Militello
    place_hemicycle: 207
    autresmandats:
      - Adjointe au Maire de Nice, Alpes-Maritimes (342482 habitants)
    mails:
      - mmarland@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267903.asp
    site_web: http://marland-militello.fr
    debut_mandat: 20/06/2007
    nom: Muriel Marland-Militello
    type: depute
  depute_267907:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 267907
    adresses:
      - Hôtel de Ville Rue de la Crouzette CS 40013 34173 Castelnau-le-Lez cedex Téléphone : 04 67 14 27 14 Télécopie : 04 67 14 27 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 34 Télécopie : 01 40 63 54 87 
      - Secrétariat parlementaire 1 Place Mendès France 34170 Castelnau-le-Lez Téléphone : 04 67 52 20 73 Télécopie : 04 67 52 29 42 
    circonscription: Hérault (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Grand
    place_hemicycle: 75
    autresmandats:
      - Membre de la communauté d'agglomération de Montpellier
      - Maire de Castelnau-le-Lez, Hérault (14214 habitants)
    mails:
      - jpgrand@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267907.asp
    profession: Attaché parlementaire
    site_web: http://www.jpgrand.com
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Grand
    type: depute
  depute_267923:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 267923
    adresses:
      - Permanence parlementaire Hôtel de ville 62307 Lens cedex Téléphone : 03 21 70 89 51 Télécopie : 03 21 70 89 51 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (13ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Delcourt
    place_hemicycle: 623
    autresmandats:
      - Maire de Lens, Pas-de-Calais (36214 habitants)
    mails:
      - delcourt.guy@laposte.net
      - gdelcourt@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267923.asp
    profession: Retraité de la fonction publique territoriale
    site_web: http://www.guydelcourt.fr
    debut_mandat: 20/06/2007
    nom: Guy Delcourt
    type: depute
  depute_267950:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléante / 
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 267950
    extras:
      - conseil national des politiques de lutte contre la pauvreté et l'exclusion sociale / membre suppléante
    adresses:
      - 14 Rue Saint-Germain-l'Auxerrois 75001 Paris Téléphone : 01 42 36 04 52 Télécopie : 01 42 36 04 53 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (1ère)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Billard
    place_hemicycle: 599
    mails:
      - mbillard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267950.asp
    profession: Bibliothécaire
    site_web: http://www.martinebillard-blog.org
    debut_mandat: 20/06/2007
    nom: Martine Billard
    type: depute
  depute_267954:
    fonctions:
      - commission des affaires européennes / membre / 
      - délégation chargée des représentants d'intérêts / membre / 
      - commission des affaires sociales / membre / 
      - délégation chargée des groupes d'études et des offices parlementaires / membre / 
      - délégation chargée de l'application du statut du député / présidente / 
      - assemblée nationale / vice-présidente / 01/10/2008
    sexe: F
    id_an: 267954
    adresses:
      - Permanence 69 Rue de la Fontaine-au-Roi 75011 Paris Téléphone : 01 43 38 76 06 Télécopie : 01 43 38 76 49 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Hoffman-Rispal
    place_hemicycle: 422
    autresmandats:
      - Membre du Conseil municipal de Paris 11ème Arrondissement, Paris (149074 habitants)
    mails:
      - dhoffman@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267954.asp
    profession: Comptable
    site_web: http://www.daniele-hoffman-rispal.fr
    debut_mandat: 20/06/2007
    nom: Danièle Hoffman-Rispal
    type: depute
  depute_267965:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 267965
    extras:
      - conseil d'administration de l'agence nationale pour la cohésion sociale et l'égalité des chances / membre suppléante
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 93 23 
      - Permanence parlementaire 30  Rue Berzélius 75017 Paris Téléphone : 01 46 27 78 32 Télécopie : 01 46 27 78 32 
    circonscription: Paris (17ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lepetit
    place_hemicycle: 450
    autresmandats:
      - Adjointe au Maire de Paris, Paris (2121291 habitants)
      - Conseillère de Paris
    mails:
      - alepetit@assemblee-nationale.fr
      - annick-lepetit@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/267965.asp
    site_web: http://www.annicklepetit.fr
    debut_mandat: 20/06/2007
    nom: Annick Lepetit
    type: depute
  depute_2679:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2679
    extras:
      - commission de vérification des fonds spéciaux (art 154 de la loi de finances pour 2002 / membre titulaire
    adresses:
      - 62 Avenue de la Châtre 36000 Châteauroux Téléphone : 02 54 08 43 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 93 16 
    circonscription: Indre (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Sapin
    place_hemicycle: 506
    autresmandats:
      - Maire d'Argenton-sur-Creuse, Indre (5151 habitants)
      - Président de la Communauté de communes du Pays d'Argenton-sur-Creuse
    mails:
      - msapin.circo@orange.fr
      - msapin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2679.asp
    profession: Conseiller de tribunal administratif
    debut_mandat: 20/06/2007
    nom: Michel Sapin
    type: depute
  depute_268001:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 268001
    extras:
      - comité national de l'eau / membre titulaire
    adresses:
      - Rue Valoise 62350 Saint-Venant Téléphone : 03 21 27 53 80 Télécopie : 03 21 27 11 56 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Flajolet
    place_hemicycle: 136
    autresmandats:
      - Maire de Saint-Venant, Pas-de-Calais (3206 habitants)
      - Membre du conseil régional (Nord-Pas-de-Calais)
    mails:
      - aflajolet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268001.asp
    profession: Professeur
    site_web: http://www.andre-flajolet.net
    debut_mandat: 20/06/2007
    nom: André Flajolet
    type: depute
  depute_268011:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 268011
    adresses:
      - Permanence parlementaire 60 Route du polygone Boîte postale A 67000 Strasbourg Téléphone : 03 88 84 55 30 Télécopie : 03 88 41 06 05 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Maurer
    place_hemicycle: 58
    autresmandats:
      - Membre du conseil général (Bas-Rhin)
    mails:
      - jmaurer@assemblee-nationale.fr
      - maurer.jean-philippe@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268011.asp
    profession: Assistant parlementaire
    site_web: http://www.jpmaurer.info
    debut_mandat: 20/06/2007
    nom: Jean-Philippe Maurer
    type: depute
  depute_268019:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - commission des lois / vice-président / 
    sexe: H
    id_an: 268019
    extras:
      - comité de l'initiative française pour les récifs coralliens / membre titulaire
    adresses:
      - Permanence parlementaire 176  Avenue Jean Jaurès 93000 Bobigny Téléphone : 01 41 50 50 50 
      - Mairie Place de l'Hôtel de Ville 93700 Drancy Téléphone : 01 48 96 50 55 Télécopie : 01 48 30 00 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (5ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Lagarde
    place_hemicycle: 367
    autresmandats:
      - Maire de Drancy, Seine-Saint-Denis (62262 habitants)
    mails:
      - jclagarde@assemblee-nationale.fr
      - lagardejc@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268019.asp
    profession: Attaché de direction
    site_web: http://www.jclagarde.net
    debut_mandat: 20/06/2007
    nom: Jean-Christophe Lagarde
    type: depute
  depute_268031:
    place_hemicycle: 466
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Maire de La Trinité, Martinique (13067 habitants)
    sexe: H
    id_an: 268031
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268031.asp
    mails:
      - ljmanscour@wanadoo.fr
      - ljmanscour@assemblee-nationale.fr
    adresses:
      - Mairie 5 Avenue Casimir Branglidor 97220 La Trinité Téléphone : 05 96 58 20 12 Télécopie : 05 96 58 65 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Martinique (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur de collège
    debut_mandat: 20/06/2007
    nom_de_famille: Manscour
    nom: Louis-Joseph Manscour
    type: depute
  depute_268039:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 268039
    adresses:
      - Dothémare 97139 Les Abymes Téléphone : 05 90 20 18 31 Télécopie : 05 90 90 48 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Guadeloupe (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Jalton
    place_hemicycle: 468
    autresmandats:
      - Maire des Abymes, Guadeloupe (63054 habitants)
      - Membre du conseil général (Guadeloupe)
    mails:
      - eric.jalton@wanadoo.fr
      - ejalton@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268039.asp
    profession: Dentiste
    site_web: http://www.ericjalton.fr
    debut_mandat: 20/06/2007
    nom: Éric Jalton
    type: depute
  depute_268042:
    place_hemicycle: 127
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire du Moule, Guadeloupe (20827 habitants)
    sexe: F
    id_an: 268042
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268042.asp
    mails:
      - glouis@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 75 Télécopie : 01 40 63 79 26 
      - Mairie Rue Joffre 97160 Le Moule Téléphone : 05 90 23 09 00 Télécopie : 05 90 23 68 73 
    circonscription: Guadeloupe (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Agent de contrôle retraitée
    debut_mandat: 20/06/2007
    nom_de_famille: Louis-Carabin
    nom: Gabrielle Louis-Carabin
    type: depute
  depute_268048:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 268048
    extras:
      - comité consultatif des liaisons aériennes d'aménagement du territoire / membre titulaire
    adresses:
      - Permanence parlementaire 6 Rue Delrieu 97100 Basse-Terre Téléphone : 05 90 80 75 15 Télécopie : 05 90 80 76 34 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Guadeloupe (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Lurel
    place_hemicycle: 505
    autresmandats:
      - Président du conseil régional (Guadeloupe)
    mails:
      - vlurel@assemblee-nationale.fr
      - victorin.lurel@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268048.asp
    profession: Fonctionnaire territorial
    site_web: http://www.lurel.parti-socialiste.fr
    debut_mandat: 20/06/2007
    nom: Victorin Lurel
    type: depute
  depute_268051:
    place_hemicycle: 190
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Maire d'Orléans, Loiret (113121 habitants)
    sexe: H
    id_an: 268051
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/268051.asp
    mails:
      - sgrouard@assemblee-nationale.fr
      - sergegrouard.deputemaire45@wanadoo.fr
    adresses:
      - Permanence parlementaire 27  Rue du Colombier 45000 Orléans Téléphone : 02 38 53 51 05 Télécopie : 02 38 77 45 02 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loiret (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Administrateur civil
    debut_mandat: 20/06/2007
    nom_de_famille: Grouard
    nom: Serge Grouard
    type: depute
  depute_2685:
    fonctions:
      - commission des affaires européennes / membre / 
      - délégation chargée des activités internationales / membre / 
      - commission des affaires étrangères / membre / 
      - délégation chargée des groupes d'études et des offices parlementaires / membre / 
      - assemblée nationale / secrétaire / 01/10/2008
    sexe: F
    id_an: 2685
    adresses:
      - 18 Rue Neyron 63000 Clermont-Ferrand Téléphone : 04 73 25 61 85 Télécopie : 04 73 24 66 41 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Puy-de-Dôme (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Saugues
    place_hemicycle: 530
    autresmandats:
      - Adjointe au Maire de Clermont-Ferrand, Puy-de-Dôme (137155 habitants)
    mails:
      - osaugues@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2685.asp
    profession: Retraitée
    site_web: http://www.odile-saugues.org
    debut_mandat: 20/06/2007
    nom: Odile Saugues
    type: depute
  depute_2690:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
      - bureau du comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: H
    id_an: 2690
    extras:
      - conseil supérieur de la sûreté et de l'information nucléaires / membre titulaire
      - conseil d'orientation de la simplification administrative / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 67 01 Télécopie : 01 40 63 52 25 
      - 12 Rue Édmé Millot 21350 Vitteaux Téléphone : 03 80 33 90 90 Télécopie : 03 80 33 90 95 
    circonscription: Côte-d'Or (4ème)
    groupe:
      - nouveau centre / président
    nom_de_famille: Sauvadet
    place_hemicycle: 364
    autresmandats:
      - Président de la communauté de communes du canton de Vitteaux
      - Président du conseil général (Côte-d'Or)
      - Adjoint au Maire de Vitteaux, Côte-d'Or (1114 habitants)
    mails:
      - francois.sauvadet@wanadoo.fr
      - fsauvadet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2690.asp
    profession: Journaliste
    site_web: http://www.francois-sauvadet.net
    debut_mandat: 20/06/2007
    nom: François Sauvadet
    type: depute
  depute_2700:
    fonctions:
      - commission des finances / membre / 
      - mission d'information commune sur l'évaluation des dispositifs fiscaux d'encouragement à l'investissement locatif / membre / 
    sexe: H
    id_an: 2700
    adresses:
      - 6 Rue du Général Leclerc BP 40049 Cedex 95210 Saint-Gratien Téléphone : 01 39 64 37 85 Télécopie : 01 39 64 37 85 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Scellier
    place_hemicycle: 290
    autresmandats:
      - Membre du conseil général (Val-d'Oise)
    mails:
      - francois.scellier@valdoise.fr
      - fscellier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2700.asp
    profession: Directeur divisionnaire des impôts honoraire
    site_web: http://www.scellier.net
    debut_mandat: 20/06/2007
    nom: François Scellier
    type: depute
  depute_2707:
    place_hemicycle: 164
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires étrangères / secrétaire / 
    sexe: H
    id_an: 2707
    extras:
      - haut conseil de la coopération internationale / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2707.asp
    mails:
      - schneider.depute@wanadoo.fr
      - aschneider@assemblee-nationale.fr
    adresses:
      - Permanence 53 Route de Bischwiller BP 12 67301 Schiltigheim cedex Téléphone : 03 88 18 55 05 Télécopie : 03 88 18 55 06 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Principal de collège en retraite
    debut_mandat: 20/06/2007
    nom_de_famille: Schneider
    nom: André Schneider
    type: depute
  depute_2708:
    place_hemicycle: 25
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Châtillon, Hauts-de-Seine (28621 habitants)
    sexe: H
    id_an: 2708
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2708.asp
    mails:
      - jpschosteck@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 Rue de l'Université 75355 Paris 07 SP 
      - Mairie de Chatillon 92320 Chatillon Téléphone : 01 42 31 81 81 Télécopie : 01 46 57 84 57 
    circonscription: Hauts-de-Seine (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 04/02/2008
    nom_de_famille: Schosteck
    nom: Jean-Pierre Schosteck
    type: depute
  depute_271:
    place_hemicycle: 523
    fonctions:
      - commission des affaires étrangères / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
    autresmandats:
      - Vice-présidente du conseil régional (Provence-Alpes-Côte-d'Azur)
    sexe: F
    id_an: 271
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/271.asp
    mails:
      - permanenceparlementaire@sylvieandrieux.fr
      - sandrieux@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 1 Place Albert Durand Village de Sainte-Marthe 13014 Marseille Téléphone : 04 95 05 15 70 Télécopie : 04 91 02 83 31 
    circonscription: Bouches-du-Rhône (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre commercial d'entreprise de manutention et d'acconage
    debut_mandat: 20/06/2007
    nom_de_famille: Andrieux
    nom: Sylvie Andrieux
    type: depute
  depute_2744:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 2744
    extras:
      - comité de suivi de la loi relative aux libertés et responsabilités des universités / membre titulaire
    adresses:
      - U.M.P. permanence 2 Bis Place Robillard 89000 Auxerre Téléphone : 03 86 52 00 98 Télécopie : 03 86 51 09 88 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 95 13 Télécopie : 01 40 63 95 39 
      - Conseil régional de Bourgogne 17 Route de la Trémouille 21000 Dijon Téléphone : 03 80 30 30 05 
      - Autre téléphone : 01 40 63 95 26  jp.soisson@wanadoo.fr
    circonscription: Yonne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Soisson
    place_hemicycle: 189
    autresmandats:
      - Membre du conseil régional (Bourgogne)
    mails:
      - jpsoisson@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2744.asp
    profession: Conseiller référendaire à la Cour des comptes
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Soisson
    type: depute
  depute_2775:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2775
    extras:
      - conseil national du tourisme / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 67 86 Télécopie : 01 40 63 54 79 
      - Mairie 21200 Beaune Téléphone : 03 80 24 56 44 Télécopie : 03 80 24 57 57 
      - Permanence 6 Place Carnot 21200 Beaune Téléphone : 03 80 22 77 80 Télécopie : 03 80 22 66 67 
    circonscription: Côte-d'Or (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Suguenot
    place_hemicycle: 294
    autresmandats:
      - Maire de Beaune, Côte-d'Or (21922 habitants)
    mails:
      - asuguenot@assemblee-nationale.fr
      - alain.suguenot@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2775.asp
    profession: Avocat
    debut_mandat: 20/06/2007
    nom: Alain Suguenot
    type: depute
  depute_2791:
    place_hemicycle: 615
    fonctions:
      - commission des affaires étrangères / membre / 
      - mission d'information commune sur les prix des carburants dans les dom / vice-présidente / 
    sexe: F
    id_an: 2791
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2791.asp
    mails:
      - ctaubira@assemblee-nationale.fr
    adresses:
      - 35  Rue Schoelcher BP 803 97300 Cayenne Téléphone : 05 94 30 31 00 Télécopie : 05 94 31 84 95 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Guyane (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    site_web: http://www.christiane-taubira.net
    profession: Économiste
    debut_mandat: 20/06/2007
    nom_de_famille: Taubira
    nom: Christiane Taubira
    type: depute
  depute_2792:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2792
    extras:
      - observatoire économique de l'achat public / membre titulaire
      - comité de gestion du fonds de soutien aux hydrocarbures ou assimiles d'origine nationale / membre titulaire
    adresses:
      - 71 Rue du Maréchal Leclerc BP 17 49250 Beaufort-en-Vallée Téléphone : 02 41 80 18 32 Télécopie : 02 41 80 18 33 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Maine-et-Loire (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Taugourdeau
    place_hemicycle: 350
    autresmandats:
      - Maire de Beaufort-en-Vallée, Maine-et-Loire (5385 habitants)
    mails:
      - jctaugourdeau.depute@wanadoo.fr
      - jctaugourdeau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2792.asp
    profession: Chef d'entreprise
    site_web: http://www.jctaugourdeau.fr
    debut_mandat: 20/06/2007
    nom: Jean-Charles Taugourdeau
    type: depute
  depute_2796:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission de la défense nationale et des forces armées / président / 
    sexe: H
    id_an: 2796
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie des 9e et 10e arrondissements 150 Boulevard Paul Claudel 13009 Marseille Téléphone : 04 91 14 63 11 Télécopie : 04 91 14 63 44 
    circonscription: Bouches-du-Rhône (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Teissier
    place_hemicycle: 168
    autresmandats:
      - Membre de la communauté urbaine Marseille Provence Métropole
      - Maire de secteur de Marseille (5ème secteur), Bouches-du-Rhône (798021 habitants)
      - Membre du Conseil municipal de Marseille, Bouches-du-Rhône (798021 habitants)
    mails:
      - gteissier@assemblee-nationale.fr
      - gteissier@mairie-marseille.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2796.asp
    profession: Administrateur de biens
    site_web: http://www.guyteissier.com
    debut_mandat: 20/06/2007
    nom: Guy Teissier
    type: depute
  depute_2799:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2799
    extras:
      - conseil de surveillance de la caisse nationale d'assurance vieillesse des travailleurs salariés / membre titulaire
      - conseil d'orientation des retraites / membre titulaire
      - conseil de surveillance de l'agence centrale des organismes de sécurité sociale / membre titulaire
      - conseil de surveillance du fonds de financement de l'allocation personnalisée d'autonomie / membre titulaire
    adresses:
      - 11 Avenue de Coux 07000 Privas Téléphone : 04 75 66 76 90 Télécopie : 04 75 66 76 91 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel du département La Chaumette 07000 Privas 
    circonscription: Ardèche (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Terrasse
    place_hemicycle: 414
    autresmandats:
      - Président du conseil général (Ardèche)
    mails:
      - pterrasse@assemblee-nationale.fr
      - pascal.terrasse@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2799.asp
    profession: Directeur de maison de retraite
    site_web: http://www.pascal-terrasse.net
    debut_mandat: 20/06/2007
    nom: Pascal Terrasse
    type: depute
  depute_2801:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2801
    adresses:
      - 8 Rue Victor Hugo 69600 Oullins Téléphone : 04 78 50 50 50 Télécopie : 04 78 86 00 44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (12ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Terrot
    place_hemicycle: 108
    autresmandats:
      - Membre du Conseil municipal d'Oullins, Rhône (25183 habitants)
    mails:
      - mterrot@michel-terrot.com
      - mterrot@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2801.asp
    profession: Avocat
    site_web: http://www.michel-terrot.com
    debut_mandat: 20/06/2007
    nom: Michel Terrot
    type: depute
  depute_2811:
    place_hemicycle: 330
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 2811
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2811.asp
    mails:
      - jeanclaude-thomas@wanadoo.fr
      - jcthomas@assemblee-nationale.fr
    adresses:
      - Secrétariat 1  Rue Roger Salengro 51100 Reims Téléphone : 03 26 40 19 20 Télécopie : 03 26 47 64 23 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Marne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Docteur en chirurgie dentaire
    debut_mandat: 20/06/2007
    nom_de_famille: Thomas
    nom: Jean-Claude Thomas
    type: depute
  depute_2815:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 2815
    extras:
      - conseil national de la formation professionnelle tout au long de la vie / membre suppléant
    adresses:
      - 486 Bis Rue Paradis 13008 Marseille Téléphone : 04 91 71 45 25 Télécopie : 04 91 76 42 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Tian
    place_hemicycle: 245
    autresmandats:
      - Maire de secteur de Marseille (4ème secteur), Bouches-du-Rhône (798021 habitants)
      - Membre du Conseil municipal de Marseille, Bouches-du-Rhône (798021 habitants)
    mails:
      - dtian@assemblee-nationale.fr
      - dominique.tian@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2815.asp
    profession: Gérant de sociétés
    debut_mandat: 20/06/2007
    nom: Dominique Tian
    type: depute
  depute_2816:
    place_hemicycle: 81
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire d'arrondissement de Paris (5ème Arrondissement), Paris (58943 habitants)
      - Conseiller de Paris, Paris (2121291 habitants)
      - Conseiller de Paris
    sexe: H
    id_an: 2816
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2816.asp
    mails:
      - jtiberi@assemblee-nationale.fr
    adresses:
      - Mairie du 5ème arrondissement 21 Place du Panthéon 75005 Paris Téléphone : 01 56 81 75 05 Télécopie : 01 56 81 75 08 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 74 Télécopie : 01 40 63 95 59 
    circonscription: Paris (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Magistrat
    debut_mandat: 20/06/2007
    nom_de_famille: Tiberi
    nom: Jean Tiberi
    type: depute
  depute_2825:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 2825
    adresses:
      - 1 Rue des Douves 37250 Montbazon Téléphone : 02 47 34 84 45 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Indre-et-Loire (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Touraine
    place_hemicycle: 432
    autresmandats:
      - Vice-présidente du conseil général (Indre-et-Loire)
    mails:
      - mtouraine@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2825.asp
    profession: Conseillère d'Etat
    site_web: http://www.marisoltouraine.typepad.fr
    debut_mandat: 20/06/2007
    nom: Marisol Touraine
    type: depute
  depute_2832:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 2832
    extras:
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Permanence parlementaire 19 Place du Général Leclerc BP 15 76760 Yerville Téléphone : 02 35 56 73 06 Télécopie : 02 35 56 13 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville Place de la Haye 76760 Yerville Téléphone : 02 32 70 43 43 Télécopie : 02 32 70 43 49 
    circonscription: Seine-Maritime (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Trassy-Paillogues
    place_hemicycle: 132
    autresmandats:
      - Président de la communauté de communes Yerville-Plateau de Caux
      - Membre du conseil général (Seine-Maritime)
      - Maire d'Yerville, Seine-Maritime (2175 habitants)
    mails:
      - atrassy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2832.asp
    profession: Ingénieur
    site_web: http://www.alfredtrassypaillogues.fr
    debut_mandat: 20/06/2007
    nom: Alfred Trassy-Paillogues
    type: depute
  depute_2843:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / coprésident / 
      - commission des finances / membre / 
    sexe: H
    id_an: 2843
    extras:
      - conseil d'orientation de l'observatoire de l'emploi public / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 05 55 
      - Hôtel de Ville BP 50 91211 Draveil cedex Téléphone : 01 69 52 78 02 Télécopie : 01 69 03 49 16 
      - Permanence 16 Avenue de la Libération 91130 Ris-Orangis Téléphone : 01 69 25 88 00 Télécopie : 01 69 06 26 58 
    circonscription: Essonne (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Tron
    place_hemicycle: 273
    autresmandats:
      - Président de la communauté d'agglomération Sénart - Val de Seine
      - Maire de Draveil, Essonne (28093 habitants)
    mails:
      - gtron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2843.asp
    profession: Agent public des collectivités locales
    site_web: http://www.georgestron.fr
    debut_mandat: 20/06/2007
    nom: Georges Tron
    type: depute
  depute_2850:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 2850
    extras:
      - conseil national de la formation professionnelle tout au long de la vie / membre titulaire
      - conseil d'administration de la société nationale de programme france 3 / membre titulaire
      - comité consultatif des liaisons aériennes d'aménagement du territoire / membre titulaire
      - commission nationale des comptes de la formation professionnelle / membre titulaire
    adresses:
      - 34 Rue de la Liberté 68300 Saint-Louis 
      - Permanence 12  Croisée des Lys 68300 Saint-Louis Téléphone : 03 89 69 15 31 Télécopie : 03 89 69 00 09 
      - Hôtel de Ville 68300 Saint-Louis Téléphone : 03 89 69 52 00 Télécopie : 03 89 69 37 72 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ueberschlag
    place_hemicycle: 167
    autresmandats:
      - Vice-président de la communauté de communes des Trois Frontières (CC3F)
      - Maire de Saint-Louis, Haut-Rhin (19961 habitants)
    mails:
      - jean.ueberschlag@wanadoo.fr
      - jueberschlag@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2850.asp
    profession: Chirurgien-dentiste retraité
    site_web: http://jean.ueberschlag.over-blog.com
    debut_mandat: 20/06/2007
    nom: Jean Ueberschlag
    type: depute
  depute_2859:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2859
    extras:
      - commission nationale de contrôle des interceptions de sécurité / membre titulaire
    adresses:
      - 13 Rue Cavé 75018 Paris Téléphone : 01 42 62 87 15 Téléphone : 01 42 54 78 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (19ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Vaillant
    place_hemicycle: 427
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Maire d'arrondissement de Paris (18ème Arrondissement), Paris (184419 habitants)
      - Conseiller de Paris
    mails:
      - dvaillant@assemblee-nationale.fr
      - contact@danielvaillant.net
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2859.asp
    profession: Technicien biologiste
    site_web: http://www.danielvaillant.net
    debut_mandat: 20/06/2007
    nom: Daniel Vaillant
    type: depute
  depute_2870:
    place_hemicycle: 498
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Président du conseil général (Isère)
    sexe: H
    id_an: 2870
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2870.asp
    mails:
      - avallini@assemblee-nationale.fr
    adresses:
      - Clos des Chartreux 38210 Tullins Téléphone : 04 76 07 96 99 Télécopie : 04 76 07 96 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (9ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Vallini
    nom: André Vallini
    type: depute
  depute_2875:
    place_hemicycle: 53
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2875
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2875.asp
    mails:
      - cvanneste@assemblee-nationale.fr
      - cvanneste@hotmail.fr
    adresses:
      - 79 Rue du Brun Pain 59200 Tourcoing Téléphone : 03 20 46 42 63 Télécopie : 03 20 94 61 09 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://vanneste.over-blog.org
    profession: Professeur de philosophie
    debut_mandat: 20/06/2007
    nom_de_famille: Vanneste
    nom: Christian Vanneste
    type: depute
  depute_2876:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2876
    extras:
      - commission d'accès aux documents administratifs / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 33 01 Télécopie : 01 40 63 33 81 
      - Permanence principale 1 Rue Baugru 88200 Remiremont Téléphone : 03 29 23 97 58 Télécopie : 03 29 23 97 60 
      - Permanence secondaire 2 Rue des Déportés 88160 Le Thillot Téléphone : 03 29 25 31 80 Télécopie : 03 29 25 35 21 
    circonscription: Vosges (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Vannson
    place_hemicycle: 341
    mails:
      - fvannson@assemblee-nationale.fr
      - f.vannson@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2876.asp
    profession: Opticien
    site_web: http://www.vannson.fr
    debut_mandat: 20/06/2007
    nom: François Vannson
    type: depute
  depute_2883:
    place_hemicycle: 417
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Président du conseil régional (Provence-Alpes-Côte-d'Azur)
    sexe: H
    id_an: 2883
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2883.asp
    mails:
      - mvauzelle@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 20 Place de la République BP 196 13637 Arles cedex Téléphone : 04 90 49 67 20 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 53 16 
    circonscription: Bouches-du-Rhône (16ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Préfet
    debut_mandat: 20/06/2007
    nom_de_famille: Vauzelle
    nom: Michel Vauzelle
    type: depute
  depute_2884:
    fonctions:
      - mission d'évaluation de la loi n°2005-370 du 22 avril 2005 relative aux droits des malades et à la fin de vie / membre / 
      - commission des lois / membre / 
    sexe: H
    id_an: 2884
    extras:
      - conseil d'orientation de la simplification administrative / membre suppléant
    adresses:
      - Permanence parlementaire,  22 Ter Cours Landrivon BP 199 13528 Port-de-Bouc cedex Téléphone : 04 42 40 54 90 Télécopie : 04 42 40 54 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (13ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Vaxès
    place_hemicycle: 589
    autresmandats:
      - Membre du Conseil municipal de Port-de-Bouc, Bouches-du-Rhône (16686 habitants)
    mails:
      - vaxes.michel@orange.fr
      - mvaxes@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2884.asp
    profession: Conseiller d'orientation-psychologue
    debut_mandat: 20/06/2007
    nom: Michel Vaxès
    type: depute
  depute_288865:
    place_hemicycle: 366
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du Conseil municipal de Bailly, Yvelines (4094 habitants)
    sexe: F
    id_an: 288865
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/288865.asp
    circonscription: Yvelines (3ème)
    groupe:
      - nouveau centre / membre
    debut_mandat: 19/04/2008
    nom_de_famille: Le Moal
    nom: Colette Le Moal
    type: depute
  depute_2895:
    place_hemicycle: 353
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Maire de Guéret, Creuse (14123 habitants)
    sexe: H
    id_an: 2895
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2895.asp
    mails:
      - mvergnier@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 64 Avenue Louis Laroche 23000 Guéret Téléphone : 05 55 52 17 17 Télécopie : 05 55 41 15 82 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Creuse (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Directeur d'école retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Vergnier
    nom: Michel Vergnier
    type: depute
  depute_2904:
    place_hemicycle: 462
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Président du conseil général (Hérault)
    sexe: H
    id_an: 2904
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2904.asp
    mails:
      - a.vezinhet.depute@orange.fr
      - avezinhet@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 100 Rue Lejzer Zamenhof Le Messidor 34080 Montpellier Téléphone : 04 67 45 02 04 Télécopie : 04 67 45 05 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hérault (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Directeur de recherche (retraité)
    debut_mandat: 20/06/2007
    nom_de_famille: Vézinhet
    nom: André Vézinhet
    type: depute
  depute_2907:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 2907
    extras:
      - conseil national du tourisme / membre titulaire
    adresses:
      - Permanence parlementaire 87 Rue de la République Les Terrasses d'Engaline 83140 Six-Fours-les-Plages Téléphone : 04 94 30 57 17 Télécopie : 04 94 34 09 03 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie Place du 18 juin BP 97 83183 Six-Fours-Les-Plages Téléphone :  04 94 34 93 69 Télécopie : 04 94 25 63 77 
    circonscription: Var (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Vialatte
    place_hemicycle: 315
    autresmandats:
      - Maire de Six-Fours-les-Plages, Var (32740 habitants)
    mails:
      - jean-sebastien.vialatte@mairie-six-fours.fr
      - jsvialatte@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2907.asp
    profession: Biologiste
    debut_mandat: 20/06/2007
    nom: Jean-Sébastien Vialatte
    type: depute
  depute_2912:
    fonctions:
      - commission des lois / vice-président / 
    sexe: H
    id_an: 2912
    adresses:
      - 11 Avenue Sadi Carnot 40000 Mont-de-Marsan Téléphone : 05 58 85 20 55 Télécopie : 05 58 06 45 67 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Landes (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Vidalies
    place_hemicycle: 354
    autresmandats:
      - Membre du conseil général (Landes)
    mails:
      - avidalies@assemblee-nationale.fr
      - alain.vidalies@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2912.asp
    profession: Avocat
    site_web: http://www.alainvidalies.fr
    debut_mandat: 20/06/2007
    nom: Alain Vidalies
    type: depute
  depute_2925:
    place_hemicycle: 553
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 2925
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2925.asp
    mails:
      - jcviollet@assemblee-nationale.fr
      - jcviollet@wanadoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 13 Boulevard de Bury 16000 Angoulême Téléphone : 05 45 93 13 70 Télécopie : 05 45 93 13 71 
    circonscription: Charente (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Assistant technique des travaux publics de l'Etat
    debut_mandat: 20/06/2007
    nom_de_famille: Viollet
    nom: Jean-Claude Viollet
    type: depute
  depute_2936:
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / secrétaire / 
      - commission de la défense nationale et des forces armées / vice-président / 
    sexe: H
    id_an: 2936
    extras:
      - commission nationale de déontologie de la sécurité / membre titulaire
    adresses:
      - Association des maires de l'Ain  45 Avenue Alsace-Lorraine BP 114 01003 Bourg-en-Bresse cedex Téléphone : 04 74 32 33 03 Télécopie : 04 74 32 58 11 
      - Mairie 01750 Replonges Téléphone : 03 85 31 18 18 Télécopie : 03 85 31 12 78 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 21 Rue de la Croix-Colin BP 28 01750 Replonges Téléphone : 03 85 31 09 70 Télécopie : 03 85 31 11 19 
    circonscription: Ain (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Voisin
    place_hemicycle: 28
    autresmandats:
      - Maire de Replonges, Ain (2845 habitants)
      - Membre du conseil régional (Rhône-Alpes)
    mails:
      - mvoisin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2936.asp
    profession: Expert comptable, commissaire aux comptes et expert-judiciaire 
    site_web: http://www.michel-voisin.net
    debut_mandat: 20/06/2007
    nom: Michel Voisin
    type: depute
  depute_2937:
    fonctions:
      - commission des affaires européennes / secrétaire / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 2937
    extras:
      - commission supérieure des sites, perspectives et paysages / membre titulaire
    adresses:
      - Mairie 71850 Charnay-lès-Mâcon  Téléphone : 03 85 34 15 70 Télécopie : 03 85 34 66 85 
      - Permanence parlementaire 3 Rue Paul Gateaud 71000 MACON Téléphone : 03.85.38.01.06 Télécopie : 03.85.39.26.50 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Voisin
    place_hemicycle: 44
    autresmandats:
      - Maire de Charnay-lès-Mâcon, Saône-et-Loire (6739 habitants)
    mails:
      - gvoisin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2937.asp
    profession: Garagiste
    site_web: http://www.gerardvoisin.com
    debut_mandat: 20/06/2007
    nom: Gérard Voisin
    type: depute
  depute_2943:
    fonctions:
      - commission des lois / secrétaire / 
    sexe: H
    id_an: 2943
    adresses:
      - Permanence 10 Avenue Jean-Baptiste Clément BP 130 08500 Revin Téléphone : 03 24 40 51 51 Télécopie : 03 24 40 51 50 
      - Autre téléphone : 01 40 63 74 60  Vuilque.Philippe@wanadoo.fr
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 74 60 
    circonscription: Ardennes (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Vuilque
    place_hemicycle: 537
    autresmandats:
      - Maire de Revin, Ardennes (8961 habitants)
    mails:
      - pvuilque@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2943.asp
    profession: Directeur de clinique
    site_web: http://www.philippevuilque.fr
    debut_mandat: 20/06/2007
    nom: Philippe Vuilque
    type: depute
  depute_2952:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des lois / président / 
    sexe: H
    id_an: 2952
    extras:
      - conseil national de l'aménagement et du développement du territoire / membre titulaire
      - conférence de la ruralité / membre titulaire
      - commission nationale de présélection des pôles d'excellence rurale / membre titulaire
    adresses:
      - Permanence 11 Rue Carnot 08200 Sedan Téléphone : 03 24 27 13 37 Télécopie : 03 24 29 12 73 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ardennes (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Warsmann
    place_hemicycle: 179
    autresmandats:
      - Président de la Communauté de communes des Trois cantons de Carignan, Mouzon et Raucourt
      - Vice-président du conseil général (Ardennes)
      - Maire de Douzy, Ardennes (1515 habitants)
    mails:
      - jlwarsmann@assemblee-nationale.fr
      - jean-luc.warsmann@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2952.asp
    profession: Sans profession
    debut_mandat: 20/06/2007
    nom: Jean-Luc Warsmann
    type: depute
  depute_295:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 295
    adresses:
      - Hôtel de Ville BP 23 93290 Tremblay-en-France Téléphone : 01 49 63 71 17 Télécopie : 01 49 63 69 66 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (11ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Asensi
    place_hemicycle: 586
    autresmandats:
      - Maire de Tremblay-en-France, Seine-Saint-Denis (33885 habitants)
    mails:
      - depute.maire@ville-tremblay-en-france.fr
      - fasensi@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/295.asp
    profession: Dessinateur industriel
    site_web: http://www.francoisasensi.com
    debut_mandat: 20/06/2007
    nom: François Asensi
    type: depute
  depute_2964:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 2964
    adresses:
      - Hôtel de ville 16 Rue du général Mangin BP K1 98849 Nouméa cedex 
      - Permanence parlementaire 13 Rue de Sébastopol BP 306 98845 Nouméa cedex 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nouvelle-Calédonie (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Yanno
    place_hemicycle: 237
    autresmandats:
      - Premier adjoint de Nouméa, Nouvelle-Calédonie (91386 habitants)
    mails:
      - gyanno@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2964.asp
    profession: Commissaire aux comptes
    site_web: http://www.yanno.nc
    debut_mandat: 20/06/2007
    nom: Gaël Yanno
    type: depute
  depute_2971:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 2971
    extras:
      - conseil de surveillance de la caisse nationale des allocations familiales / membre titulaire
    circonscription: Moselle (3ème)
    adresses:
      - 9 Square du Pontiffroy 57000 Metz Téléphone : 03 87 30 39 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Zimmermann
    place_hemicycle: 36
    autresmandats:
      - Membre du conseil régional (Lorraine)
      - Membre du Conseil municipal de Metz, Moselle (123776 habitants)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/2971.asp
    mails:
    profession: Professeur certifié
    debut_mandat: 20/06/2007
    nom: Marie-Jo Zimmermann
    type: depute
  depute_303108:
    place_hemicycle: 56
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 303108
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/303108.asp
    circonscription: Haute-Loire (1ère)
    groupe:
      - union pour un mouvement populaire / apparenté
    profession: Cadre bancaire
    debut_mandat: 20/07/2007
    nom_de_famille: Marcon
    nom: Jean-Pierre Marcon
    type: depute
  depute_304016:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 304016
    adresses:
      - 42 Boulevard du Général de Gaulle 76200 Dieppe Téléphone : 02 35 06 11 52 Télécopie : 02 35 06 12 14 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 31 13 Télécopie : 01 40 63 31 93 
    circonscription: Seine-Maritime (11ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Hurel
    place_hemicycle: 633
    autresmandats:
      - Membre du conseil général (Seine-Maritime)
    mails:
      - sandrine.hurel@cg76.fr
      - hurel.sandrine@wanadoo.fr
      - shurel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/304016.asp
    profession: Secrétaire de direction
    site_web: http://sandrine-hurel.info
    debut_mandat: 20/06/2007
    nom: Sandrine Hurel
    type: depute
  depute_309643:
    place_hemicycle: 66
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Vice-présidente du conseil général (Vendée)
    sexe: F
    id_an: 309643
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/309643.asp
    mails:
      - vbesse@assemblee-nationale.fr
      - veronique.besse@vendee.fr
    adresses:
      - 14  Rue de Saumur 85500 Les Herbiers Téléphone : 02 51 92 94 95 Télécopie : 02 51 92 94 96 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vendée (4ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Besse
    nom: Véronique Besse
    type: depute
  depute_312:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 312
    adresses:
      - Mairie 23140 Cressat Téléphone : 05 55 62 93 59 Télécopie : 05 55 62 33 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Creuse (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Auclair
    place_hemicycle: 60
    autresmandats:
      - Maire de Cressat, Creuse (523 habitants)
      - Membre du conseil général (Creuse)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/312.asp
    mails:
      - auclair.j@wanadoo.fr
    site_web: http://www.jean-auclair.fr
    profession: Agriculteur
    debut_mandat: 20/06/2007
    nom: Jean Auclair
    type: depute
  depute_320:
    fonctions:
      - commission des affaires étrangères / vice-présidente / 
    sexe: F
    id_an: 320
    extras:
      - conseil supérieur de la coopération / membre titulaire
      - conseil d'administration de l'etablissement public du musée du quai branly / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Aurillac
    place_hemicycle: 182
    mails:
      - maurillac@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/320.asp
    profession: Attachée d'administration centrale en détachement
    site_web: http://www.martine-aurillac.fr
    debut_mandat: 20/06/2007
    nom: Martine Aurillac
    type: depute
  depute_328:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
      - bureau du comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: H
    id_an: 328
    extras:
      - comité d'orientation du centre d'analyse stratégique / membre titulaire
    adresses:
      - Permanence parlementaire 47  Place de Preux BP 351 44816 Saint-Herblain Cedex Téléphone : 02 40 43 13 18 Télécopie : 02 40 46 15 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / président
    nom_de_famille: Ayrault
    place_hemicycle: 508
    autresmandats:
      - Président de la communauté urbaine de Nantes Métropole
      - Maire de Nantes, Loire-Atlantique (269131 habitants)
    mails:
      - jmayrault@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/328.asp
    profession: Professeur d'allemand
    debut_mandat: 20/06/2007
    nom: Jean-Marc Ayrault
    type: depute
  depute_330008:
    place_hemicycle: 50
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du Conseil municipal de Bourg-en-Bresse, Ain (40666 habitants)
    sexe: H
    id_an: 330008
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330008.asp
    mails:
      - contact@xavier-breton.com
      - xbreton@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 27 Rue du Docteur Hudellet 01000 Bourg-en-Bresse Téléphone : 04 74 45 02 11 Télécopie : 04 74 22 37 07 
    circonscription: Ain (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre territorial
    debut_mandat: 20/06/2007
    nom_de_famille: Breton
    nom: Xavier Breton
    type: depute
  depute_330112:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 330112
    adresses:
      - Permanence parlementaire 6 Bis  rue du général de Gaulle 02400 Château-Thierry 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aisne (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Vasseur
    place_hemicycle: 236
    autresmandats:
      - Vice-présidente Union des communautés de communes du sud de l'Aisne
      - Maire de Ronchères, Aisne (121 habitants)
      - Membre du conseil général (Aisne)
    mails:
      - ivasseur@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330112.asp
    profession: Infirmière
    site_web: http://www.isabellevasseur.fr
    debut_mandat: 20/06/2007
    nom: Isabelle Vasseur
    type: depute
  depute_330118:
    place_hemicycle: 650
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire d'Yzeure, Allier (12696 habitants)
      - Vice-président de Moulins Communauté
    sexe: H
    id_an: 330118
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330118.asp
    mails:
      - guy.chambefort@orange.fr
      - gchambefort@assemblee-nationale.fr
    adresses:
      - Mairie d'Yzeure Place Jules Ferry 03400 Yzeure Téléphone : 04 70 20 23 68 Télécopie : 04 70 46 10 81 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Allier (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    profession: Retraité de l'enseignement
    debut_mandat: 20/06/2007
    nom_de_famille: Chambefort
    nom: Guy Chambefort
    type: depute
  depute_330130:
    place_hemicycle: 487
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 330130
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330130.asp
    mails:
      - bernard.lesterlin@orange.fr
      - blesterlin@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 148 Bis Boulevard de Courtais 03100 Montluçon Téléphone : 04 70 03 74 31 Télécopie : 04 70 09 31 22 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Allier (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://bernardlesterlin.typepad.fr
    profession: Administrateur civil
    debut_mandat: 20/06/2007
    nom_de_famille: Lesterlin
    nom: Bernard Lesterlin
    type: depute
  depute_330146:
    fonctions:
      - commission des affaires sociales / secrétaire / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / coprésident / 
      - comité d'évaluation et de contrôle des politiques publiques / vice-président / 
    sexe: H
    id_an: 330146
    adresses:
      - Permanence parlementaire 60 Rue Victor Hugo 03500 Saint-Pourçain-sur-Sioule Téléphone : 04 70 45 44 68 Télécopie : 04 70 47 53 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Allier (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Mallot
    place_hemicycle: 488
    autresmandats:
      - Membre du conseil régional (Auvergne)
    mails:
      - jmallot@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330146.asp
    profession: Contrôleur général économique et financier
    site_web: http://jean.mallot.over-blog.com
    debut_mandat: 20/06/2007
    nom: Jean Mallot
    type: depute
  depute_330240:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 330240
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 96 Télécopie : 01 40 63 78 41 
      - 13 Rue Saint François de Paule 06300 Nice Téléphone : 04 93 85 22 26 Télécopie : 04 93 85 20 79 
    circonscription: Alpes-Maritimes (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Ciotti
    place_hemicycle: 155
    autresmandats:
      - Président du conseil général (Alpes-Maritimes)
    mails:
      - e.ciotti@orange.fr
      - eciotti@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330240.asp
    profession: Directeur de cabinet d'un président de conseil général
    site_web: http://www.eric-ciotti.fr
    debut_mandat: 20/06/2007
    nom: Éric Ciotti
    type: depute
  depute_330357:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 330357
    adresses:
      - 1 Rue Sadi Carnot 07100 Annonay 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ardèche (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Dussopt
    place_hemicycle: 381
    autresmandats:
      - Maire d'Annonay, Ardèche (17522 habitants)
    mails:
      - odussopt@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330357.asp
    profession: Assistant parlementaire
    site_web: http://www.olivierdussopt.fr
    debut_mandat: 20/06/2007
    nom: Olivier Dussopt
    type: depute
  depute_330546:
    place_hemicycle: 570
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Membre du conseil régional (Midi-Pyrénées)
    sexe: F
    id_an: 330546
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330546.asp
    mails:
      - mlmarcel@assemblee-nationale.fr
      - marielou.marcel.p@orange.fr
    adresses:
      - 6 Avenue du Quercy 12200 Villefranche de Rouergue Téléphone : 05 65 45 62 25 
      - 20 Rue Emma Calvé 12300 Decazeville Téléphone : 05 65 43 02 27 Télécopie : 05 65 63 92 24 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aveyron (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Responsable Ressources Humaines en dispense d'activité
    debut_mandat: 20/06/2007
    nom_de_famille: Marcel
    nom: Marie-Lou Marcel
    type: depute
  depute_330613:
    fonctions:
      - commission des affaires économiques / membre / 
      - mission d'information commune sur l'indemnisation des victimes des maladies nosocomiales et accès au dossier médical / membre / 
    sexe: H
    id_an: 330613
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Conseil général des Bouches du Rhône 52 Avenue de Saint Just 13004 Marseille 
    circonscription: Bouches-du-Rhône (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Jibrayel
    place_hemicycle: 394
    autresmandats:
      - Membre du conseil général (Bouches-du-Rhône)
    mails:
      - hjibrayel@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330613.asp
    profession: Retraité des entreprises publiques
    site_web: http://henrijibrayel.over-blog.com
    debut_mandat: 20/06/2007
    nom: Henri Jibrayel
    type: depute
  depute_330684:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 330684
    extras:
      - conseil de surveillance du fonds de réserve pour les retraites / membre suppléante
    adresses:
      - 99 Avenue de la Rose 13013 Marseille Téléphone : 04 91 06 54 33 Télécopie : 04 91 06 54 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Boyer
    place_hemicycle: 223
    autresmandats:
      - Adjointe au Maire de Marseille, Bouches-du-Rhône (798021 habitants)
    mails:
      - vboyer@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330684.asp
    profession: Cadre du secteur hospitalier
    site_web: http://www.valerieboyer.fr
    debut_mandat: 20/06/2007
    nom: Valérie Boyer
    type: depute
  depute_330788:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 330788
    extras:
      - conseil stratégique du commerce de proximité / membre titulaire
    adresses:
      - 34 Avenue du général de Gaulle 13160 Châteaurenard Téléphone : 04.32.62.10.06 Télécopie : 04.32.61.08.44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (15ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Reynès
    place_hemicycle: 12
    autresmandats:
      - Vice-président Communauté de communes Rhône - Alpilles - Durance
      - Maire de Châteaurenard, Bouches-du-Rhône (13070 habitants)
    mails:
      - breynes@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330788.asp
    profession: Dentiste
    site_web: http://www.bernard-reynes.com
    debut_mandat: 20/06/2007
    nom: Bernard Reynès
    type: depute
  depute_330909:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 330909
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 21 Rue des Frères 15000 Aurillac Téléphone : 04 71 43 31 00 Télécopie : 04 71 43 13 00 
    circonscription: Cantal (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Descoeur
    place_hemicycle: 49
    autresmandats:
      - Président du conseil général (Cantal)
      - Membre du Conseil municipal de Montsalvy, Cantal (896 habitants)
    mails:
      - vdescoeur@cg15.fr
      - vdescoeur@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330909.asp
    profession: Professeur agrégé de biologie
    site_web: http://www.descoeur.com
    debut_mandat: 20/06/2007
    nom: Vincent Descoeur
    type: depute
  depute_330981:
    place_hemicycle: 649
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Adjointe au Maire de Balzac, Charente (1237 habitants)
    sexe: F
    id_an: 330981
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/330981.asp
    mails:
      - mpinville@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 7 Place de l'Hôtel de ville 16160 Gond Pontouvre Téléphone : 05 45 90 33 90 Télécopie : 05 45 95 86 59 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Charente (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    profession: Retraitée de la fonction publique
    debut_mandat: 20/06/2007
    nom_de_famille: Pinville
    nom: Martine Pinville
    type: depute
  depute_331014:
    place_hemicycle: 482
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / secrétaire / 
    sexe: F
    id_an: 331014
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331014.asp
    mails:
      - cquere@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 2 Rue René Cassin 17100 Saintes Téléphone : 05 46 91 69 42 Télécopie : 05 46 92 97 16 
      - 8 Boulevard Jacques Caillaud 17400 Saint Jean d'Angely 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 62 59 
    circonscription: Charente-Maritime (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.catherine-quere.fr
    profession:  Viticultrice
    debut_mandat: 20/06/2007
    nom_de_famille: Catherine Quéré
    nom: Catherine Quéré
    type: depute
  depute_331146:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 331146
    adresses:
      - Hôtel de ville,  20620 Biguglia Téléphone : 04 95 58 98 58 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Corse (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gandolfi-Scheit
    place_hemicycle: 244
    autresmandats:
      - Maire de Biguglia, Haute-Corse (6200 habitants)
    mails:
      - sgandolfi@assemblee-nationale.fr
      - depute-gandolfi@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331146.asp
    profession: Médecin
    site_web: http://www.depute-gandolfi.com
    debut_mandat: 20/06/2007
    nom: Sauveur Gandolfi-Scheit
    type: depute
  depute_331282:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 331282
    adresses:
      - Résidence du Manoir 32 Bis Place du Marchallac'h 22300 Lannion Téléphone : 02 96 37 03 23 Télécopie : 02 96 37 05 70 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côtes-d'Armor (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Erhel
    place_hemicycle: 565
    autresmandats:
      - Membre du conseil régional (Bretagne)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331282.asp
    mails:
      - erhel.corinne@orange.fr
    site_web: http://www.corinne-erhel.fr
    profession: Assistante parlementaire
    debut_mandat: 20/06/2007
    nom: Corinne Erhel
    type: depute
  depute_331381:
    place_hemicycle: 48
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 331381
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331381.asp
    mails:
      - jgrosperrin@assemblee-nationale.fr
    adresses:
      - Permanence 9 Avenue Edouard Droz 25000 Besançon Téléphone : 03 81 51 98 88 Télécopie : 03 81 52 13 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Doubs (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.grosperrin.net
    profession: Professeur de faculté
    debut_mandat: 20/06/2007
    nom_de_famille: Grosperrin
    nom: Jacques Grosperrin
    type: depute
  depute_331442:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 331442
    adresses:
      - Hôtel de ville Place Emile Loubet 26200 Montélimar Téléphone : 04 75 00 25 05 Télécopie : 04 75 00 25 72 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Drôme (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Reynier
    place_hemicycle: 241
    autresmandats:
      - Maire de Montélimar, Drôme (31344 habitants)
      - Président de la Communauté de communes de l'Agglomération de Montélimar
    mails:
      - freynier@assemblee-nationale.fr
      - courriel@franck-reynier.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331442.asp
    profession: Informaticien
    site_web: http://www.franck-reynier.fr
    debut_mandat: 20/06/2007
    nom: Franck Reynier
    type: depute
  depute_331567:
    fonctions:
      - commission des affaires économiques / vice-présidente / 
    sexe: F
    id_an: 331567
    extras:
      - commission du dividende numérique / membre titulaire
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Permanence 6 Allée Édouard Manet 28110 Lucé Téléphone : 02 37 34 84 29 Télécopie : 02 37 28 24 02 
      - Permanence 17 Clos Couronnet 28400 Nogent-le-Rotrou Téléphone : 02 37 52 10 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 72 53 
    circonscription: Eure-et-Loir (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Laure de La Raudière
    place_hemicycle: 322
    autresmandats:
      - Vice-présidente de la communauté de communes du Pays Courvillois
      - Adjointe au Maire de Saint-Denis-des-Puits, Eure-et-Loir (116 habitants)
    mails:
      - ldelaraudiere@assemblee-nationale.fr
      - laure@la-raudiere.com
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331567.asp
    profession: Chef d'entreprise
    site_web: http://www.la-raudiere.com
    debut_mandat: 20/06/2007
    nom: Laure de La Raudière
    type: depute
  depute_331582:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 331582
    adresses:
      - Permanence parlementaire Rue André Gillet 28200 Châteaudun Téléphone : 02 37 45 28 24 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Eure-et-Loir (4ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Vigier
    place_hemicycle: 388
    autresmandats:
      - Maire de Cloyes-sur-le-Loir, Eure-et-Loir (2645 habitants)
      - Membre du conseil régional (Centre)
    mails:
      - pvigier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331582.asp
    profession: Médecin
    site_web: http://www.philippevigier.com
    debut_mandat: 20/06/2007
    nom: Philippe Vigier
    type: depute
  depute_331594:
    place_hemicycle: 486
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission des lois / membre / 
    sexe: H
    id_an: 331594
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331594.asp
    mails:
      - contact@urvoas.org
      - jjurvoas@assemblee-nationale.fr
    adresses:
      - 8-10 Place de la Tourbie 29000 Quimper Téléphone : 02 98 95 69 80 Télécopie : 02 98 95 01 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Finistère (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.urvoas.org
    profession: Maître de conférences
    debut_mandat: 20/06/2007
    nom_de_famille: Urvoas
    nom: Jean-Jacques Urvoas
    type: depute
  depute_331658:
    fonctions:
      - commission des affaires économiques / secrétaire / 
    sexe: F
    id_an: 331658
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 12 Rue du Prat Résidence Pierre Pichavant 29120 Pont-l'Abbé Téléphone : 02 98 82 31 68 Télécopie : 02 98 87 31 08 
    circonscription: Finistère (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Loch
    place_hemicycle: 485
    autresmandats:
      - Membre du conseil général (Finistère)
    mails:
      - annick.leloch.deputee@orange.fr
      - aleloch@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331658.asp
    profession: Commercant
    site_web: http://www.annickleloch.fr
    debut_mandat: 20/06/2007
    nom: Annick Le Loch
    type: depute
  depute_331753:
    place_hemicycle: 572
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 331753
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331753.asp
    mails:
      - catherine.lemorton@orange.fr
      - clemorton@assemblee-nationale.fr
    adresses:
      - 47 Bis Boulevard de Strasbourg 31000 Toulouse Téléphone : 05 61 13 76 50 Télécopie : 05 61 12 44 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://catherine-lemorton.eu
    profession: Pharmacien
    debut_mandat: 20/06/2007
    nom_de_famille: Lemorton
    nom: Catherine Lemorton
    type: depute
  depute_331807:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 331807
    adresses:
      - Permanence parlementaire 37 Rue Clément Ader 31300 Toulouse Téléphone : 05 34 26 51 85 Télécopie : 05 34 26 13 42 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Martinel
    place_hemicycle: 571
    autresmandats:
      - Membre du conseil général (Haute-Garonne)
    mails:
      - mmartinel@assemblee-nationale.fr
      - martinemartinel@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331807.asp
    profession: Enseignant
    site_web: http://www.martine-martinel.org
    debut_mandat: 20/06/2007
    nom: Martine Martinel
    type: depute
  depute_331835:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 331835
    adresses:
      - 50 Avenue Marie Curie 31600 Seysses Téléphone : 05 61 44 63 82 Télécopie : 05 61 08 84 68 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Iborra
    place_hemicycle: 463
    autresmandats:
      - Premier Vice-président du conseil régional (Midi-Pyrénées)
    mails:
      - miborra@assemblee-nationale.fr
      - monique.iborra@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331835.asp
    profession: Fonctionnaire de catégorie A
    site_web: http://www.moniqueiborra.net
    debut_mandat: 20/06/2007
    nom: Monique Iborra
    type: depute
  depute_331924:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 331924
    adresses:
      - Permanence parlementaire 20 Rue Saint Laurent 33000 Bordeaux Téléphone : 05 56 44 84 80 Télécopie : 05 56 52 57 06 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Delaunay
    place_hemicycle: 383
    autresmandats:
      - Membre du conseil général (Gironde)
    mails:
      - delaunay.deputee@orange.fr
      - mdelaunay@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331924.asp
    profession: Médecin des hôpitaux
    site_web: http://www.michele-delaunay.net
    debut_mandat: 20/06/2007
    nom: Michèle Delaunay
    type: depute
  depute_331973:
    place_hemicycle: 382
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 331973
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331973.asp
    mails:
      - pgot@assemblee-nationale.fr
      - contact@pascalegot.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 03 13 
      - Bureau de poste principal BP 30 33320 Eysines Téléphone : 05 56 15 65 28 Télécopie : 05 56 15 51 36 
    circonscription: Gironde (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.pascalegot.fr
    profession: Journaliste
    debut_mandat: 20/06/2007
    nom_de_famille: Got
    nom: Pascale Got
    type: depute
  depute_331990:
    place_hemicycle: 418
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Président du conseil régional (Aquitaine)
    sexe: H
    id_an: 331990
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/331990.asp
    mails:
      - arousset@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 00 Télécopie : 01 40 63 93 93 
      - Permanence Hôtel de ville Place de la Ve République 33604 PESSAC cedex Téléphone : 09 62 26 14 03 
    circonscription: Gironde (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre supérieur (secteur privé)
    debut_mandat: 20/06/2007
    nom_de_famille: Rousset
    nom: Alain Rousset
    type: depute
  depute_332015:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 332015
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (9ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Faure
    place_hemicycle: 642
    autresmandats:
      - Membre du Conseil municipal d'Aillas, Gironde (668 habitants)
      - Membre du conseil général (Gironde)
    mails:
      - martine.faure2007@orange.fr
      - mfaure@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332015.asp
    profession: Retraitée de l'enseignement
    site_web: http://www.martinefaure.fr
    debut_mandat: 20/06/2007
    nom: Martine Faure
    type: depute
  depute_332154:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 332154
    extras:
      - commission supérieure du crédit maritime mutuel / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Hérault (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: d'Ettore
    place_hemicycle: 124
    autresmandats:
      - Maire d'Agde, Hérault (19988 habitants)
      - Président de la communauté d'agglomération Hérault Méditerranée
    mails:
      - gdettore@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332154.asp
    profession: Permanent politique
    site_web: http://www.gillesdettore.fr
    debut_mandat: 20/06/2007
    nom: Gilles d'Ettore
    type: depute
  depute_332206:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 332206
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 55 Rue Notre Dame 35600 Redon 
    circonscription: Ille-et-Vilaine (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Marsac
    place_hemicycle: 484
    autresmandats:
      - Membre du conseil régional (Bretagne)
    mails:
      - jrmarsac@assemblee-nationale.fr
      - jrmarsac.permanence@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332206.asp
    profession: Cadre
    site_web: http://www.jrmarsac-leblog.typepad.fr
    debut_mandat: 20/06/2007
    nom: Jean-René Marsac
    type: depute
  depute_332228:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 332228
    adresses:
      - 1 Bis Boulevard Leclerc 35300 Fougères Téléphone : 02 99 17 11 71 Télécopie : 02 99 17 11 72 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ille-et-Vilaine (6ème)
    groupe:
      - nouveau centre / apparenté
    nom_de_famille: Benoit
    place_hemicycle: 402
    autresmandats:
      - Adjoint au Maire de Lécousse, Ille-et-Vilaine (2821 habitants)
    mails:
      - thierry.benoit13@wanadoo.fr
      - tbenoit@assemblee-nationale.fr
      - contact@thierry-benoit.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332228.asp
    profession: Représentant de commerce
    site_web: http://www.thierry-benoit.fr
    debut_mandat: 20/06/2007
    nom: Thierry Benoit
    type: depute
  depute_332305:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 332305
    extras:
      - conseil national de la formation professionnelle tout au long de la vie / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 69 49 
      - Permanence parlementaire 45 Avenue de Grammont 37000 Tours Téléphone : 02 47 20 25 28 Télécopie : 02 47 20 25 29 
    circonscription: Indre-et-Loire (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Gille
    place_hemicycle: 395
    autresmandats:
      - Membre du Conseil municipal de Tours, Indre-et-Loire (132820 habitants)
    mails:
      - jpgille@assemblee-nationale.fr
      - contact@jean-patrick-gille.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332305.asp
    profession: Chargé de mission auprès d'un conseil régional
    site_web: http://blog.jean-patrick-gille.fr/
    debut_mandat: 20/06/2007
    nom: Jean-Patrick Gille
    type: depute
  depute_332364:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 332364
    extras:
      - conseil d'administration de l'agence nationale pour la gestion des déchets radioactifs / membre titulaire
    adresses:
      - Permanence 7 Rue Voltaire 38000 Grenoble 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Fioraso
    place_hemicycle: 568
    autresmandats:
      - Adjointe au Maire de Grenoble, Isère (153298 habitants)
      - Vice-présidente de la communauté d'agglomération Grenoble-Alpes Métropole
    mails:
      - genevieve.fioraso@gmail.com
      - gfioraso@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332364.asp
    profession: Cadre supérieur
    site_web: http://www.genevieve-fioraso.fr
    debut_mandat: 20/06/2007
    nom: Geneviève Fioraso
    type: depute
  depute_332384:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'information commune sur les exonérations sociales / membre / 
    sexe: H
    id_an: 332384
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 21 Rue du Doyen Gosse 38400 Saint Martin d'Hères Téléphone : 04 76 57 04 37 Télécopie : 04 76 41 84 04 
    circonscription: Isère (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Issindou
    place_hemicycle: 483
    autresmandats:
      - Maire de Gières, Isère (6232 habitants)
      - Vice-président de la communauté d'agglomération Grenoble-Alpes Métropole
    mails:
      - missindou@assemblee-nationale.fr
      - michel.issindou@free.fr
      - michel.issindou@ville-gieres.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332384.asp
    profession: Cadre de la fonction publique
    site_web: http://issindou.unblog.fr
    debut_mandat: 20/06/2007
    nom: Michel Issindou
    type: depute
  depute_332523:
    place_hemicycle: 39
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Membre du conseil général (Jura)
    sexe: F
    id_an: 332523
    extras:
      - conseil supérieur de la forêt, des produits forestiers et de la transformation du bois / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332523.asp
    mails:
      - marie-christine.dalloz390@orange.fr
      - mcdalloz@assemblee-nationale.fr
      - marie-christine.dalloz39@orange.fr
    adresses:
      - 63 Rue du Collège 39200 Saint-Claude Téléphone : 03 84 45 11 14 
      - 2 Rue du Général Leclerc 39300 Champagnole Téléphone : 03 84 52 05 13 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Jura (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Dalloz
    nom: Marie-Christine Dalloz
    type: depute
  depute_332614:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 332614
    adresses:
      - 11 Rue de la Résistance 42000 Saint-Etienne Téléphone : 04 77 30 53 60 Télécopie : 04 77 30 94 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 15 62 Télécopie : 01 40 63 15 64 
    circonscription: Loire (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Juanico
    place_hemicycle: 564
    autresmandats:
      - Membre du conseil général (Loire)
    mails:
      - rjuanico@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332614.asp
    profession: Fonctionnaire territorial
    site_web: http://www.juanico.fr
    debut_mandat: 20/06/2007
    nom: Régis Juanico
    type: depute
  depute_332636:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / membre / 
      - commission des affaires économiques / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
    sexe: H
    id_an: 332636
    adresses:
      - 2 Rue Faure-Belon BP 60 208 42005 Saint-Étienne cedex 1 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Gagnaire
    place_hemicycle: 393
    autresmandats:
      - Vice-président du conseil régional (Rhône-Alpes)
    mails:
      - contact@jlgagnaire.com
      - jlgagnaire@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332636.asp
    profession: Enseignant
    site_web: http://www.jlgagnaire.com
    debut_mandat: 20/06/2007
    nom: Jean-Louis Gagnaire
    type: depute
  depute_332747:
    fonctions:
      - assemblée nationale / secrétaire / 27/06/2007
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - comité d'évaluation et de contrôle des politiques publiques / secrétaire / 
      - commission des finances / membre / 
      - délégation chargée de l'application du statut du député / membre / 
    sexe: H
    id_an: 332747
    extras:
      - commission nationale pour l'autonomie des jeunes / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 90 Rue Paul Bellamy 44000 Nantes 
    circonscription: Loire-Atlantique (1ère)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Rugy
    place_hemicycle: 601
    autresmandats:
      - Membre du Conseil municipal d'Orvault, Loire-Atlantique (23558 habitants)
      - Membre de la communauté urbaine de Nantes Métropole
    mails:
      - permanence.fderugy@orange.fr
      - fderugy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332747.asp
    profession: Assistant parlementaire
    site_web: http://blog.francoisderugy.fr
    debut_mandat: 20/06/2007
    nom: François de Rugy
    type: depute
  depute_332796:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / membre / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 332796
    adresses:
      - Permanence parlementaire 4 Rue Léonard de Vinci 44470 Carquefou 
    circonscription: Loire-Atlantique (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Ménard
    place_hemicycle: 604
    autresmandats:
      - Membre du conseil général (Loire-Atlantique)
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332796.asp
    mails:
      - contact@michelmenard.fr
    site_web: http://www.michelmenard.fr
    profession: Professeur des écoles
    debut_mandat: 20/06/2007
    nom: Michel Ménard
    type: depute
  depute_332843:
    place_hemicycle: 603
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Vice-présidente de la communauté d'agglomération de la région nazairienne et l'estuaire
      - Membre du Conseil municipal de Saint-Nazaire, Loire-Atlantique (65874 habitants)
    sexe: F
    id_an: 332843
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332843.asp
    mails:
      - mobouille@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 30 Rue de Bois Savary BP 50132 44603 Saint-Nazaire Cedex Téléphone : 02 51 10 10 51 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Sage-femme
    debut_mandat: 20/06/2007
    nom_de_famille: Marie-Odile Bouillé
    nom: Marie-Odile Bouillé
    type: depute
  depute_332858:
    place_hemicycle: 319
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    autresmandats:
      - Maire de Pornic, Loire-Atlantique (11899 habitants)
    sexe: H
    id_an: 332858
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332858.asp
    mails:
      - pboennec@assemblee-nationale.fr
    adresses:
      - 12, Rue Sainte-Victoire 44210 Pornic Téléphone : 02 28 53 04 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin
    debut_mandat: 20/06/2007
    nom_de_famille: Boënnec
    nom: Philippe Boënnec
    type: depute
  depute_332886:
    place_hemicycle: 63
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / membre / 
      - commission des affaires économiques / membre / 
    autresmandats:
      - Premier adjoint d'Orléans, Loiret (113121 habitants)
    sexe: H
    id_an: 332886
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332886.asp
    mails:
      - ocarre@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 491 Rue Marcel Belot 45160 Olivet Téléphone : 02 38 69 03 07 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loiret (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chef d'entreprise
    debut_mandat: 20/06/2007
    nom_de_famille: Olivier Carré
    nom: Olivier Carré
    type: depute
  depute_332950:
    place_hemicycle: 630
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Membre du conseil général (Lot)
    sexe: F
    id_an: 332950
    mails:
      - orliacdominique@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/332950.asp
    circonscription: Lot (1ère)
    adresses:
      - Permanence parlementaire 93 Rue Caviole BP 233 46000 Cahors Téléphone : 05 65 35 01 08 Télécopie : 05 65 35 04 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    profession: Médecin
    debut_mandat: 20/06/2007
    nom_de_famille: Orliac
    nom: Dominique Orliac
    type: depute
  depute_333043:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 333043
    adresses:
      - Hôtel de ville BP 27 49800 Trélazé Téléphone : 02 41 33 74 60 Télécopie : 02 41 69 71 73 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Maine-et-Loire (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Goua
    place_hemicycle: 406
    autresmandats:
      - Maire de Trélazé, Maine-et-Loire (11016 habitants)
    mails:
      - secretariat.mairie@mairie-trelaze.fr
      - mgoua@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333043.asp
    profession: Retraité salarié privé
    site_web: http://www.marcgoua.fr
    debut_mandat: 20/06/2007
    nom: Marc Goua
    type: depute
  depute_333134:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - mission d'information commune sur l'indemnisation des victimes des maladies nosocomiales et accès au dossier médical / président / 
      - commission des lois / membre / 
    sexe: H
    id_an: 333134
    adresses:
      - 22 Rue du Jardin des Plantes 50300 Avranches Téléphone : 02 33 60 99 38 Télécopie : 02 33 48 75 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie Place Littré 50300 Avranches Téléphone : 02 33 89 29 52 Télécopie : 02 33 58 17 90 
    circonscription: Manche (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Huet
    place_hemicycle: 149
    autresmandats:
      - Maire d'Avranches, Manche (8500 habitants)
      - Président de la communauté de communes du canton d'Avranches
    mails:
      - ghuet@assemblee-nationale.fr
      - guenhael.huet@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333134.asp
    profession: Fonctionnaire
    site_web: http://www.guenael-huet.org
    debut_mandat: 20/06/2007
    nom: Guénhaël Huet
    type: depute
  depute_333224:
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Adjoint au Maire de Châlons-en-Champagne, Marne (47339 habitants)
    sexe: H
    id_an: 333224
    extras:
      - comité de suivi de la loi relative aux libertés et responsabilités des universités / membre suppléant
      - conseil d'administration du centre national des oeuvres universitaires et scolaires / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333224.asp
    mails:
      - bapparu@assemblee-nationale.fr
      - contact@benoistapparu.com
    adresses:
      - Permanence parlementaire 25 Rue Prieur de la Marne 51000 Châlons-en-Champagne Téléphone : 03 26 64 13 12 Télécopie : 03 26 64 79 79 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Marne (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.benoistapparu.com
    debut_mandat: 20/06/2007
    nom_de_famille: Apparu
    nom: Benoist Apparu
    type: depute
  depute_333285:
    place_hemicycle: 566
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Laval, Mayenne (50947 habitants)
      - Président de la communauté d'agglomération de Laval
    sexe: H
    id_an: 333285
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333285.asp
    mails:
      - ggarot@assemblee-nationale.fr
    adresses:
      - 22 Rue Souchu-Servinière 53000 Laval Téléphone : 02 43 01 03 05 Télécopie : 02 43 01 17 10 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Mayenne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Garot
    nom: Guillaume Garot
    type: depute
  depute_333335:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 333335
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meurthe-et-Moselle (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Féron
    place_hemicycle: 645
    autresmandats:
      - Maire de Tomblaine, Meurthe-et-Moselle (7853 habitants)
    mails:
      - hferon@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333335.asp
    profession: Homme de lettres et Artiste
    site_web: http://herveferon.fr
    debut_mandat: 20/06/2007
    nom: Hervé Féron
    type: depute
  depute_333352:
    place_hemicycle: 144
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires sociales / membre / 
    autresmandats:
      - Adjointe au Maire de Nancy, Meurthe-et-Moselle (103606 habitants)
      - Membre de la communauté urbaine du Grand Nancy
    sexe: F
    id_an: 333352
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333352.asp
    mails:
      - permanence@v-r-d.fr
      - vrosso@assemblee-nationale.fr
    adresses:
      - 23 Rue Lavigerie Bâtiment B 54000 Nancy Téléphone : 03 83 41 69 20 Télécopie : 03 83 41 12 98 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Meurthe-et-Moselle (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Juriste d'entreprise
    debut_mandat: 20/06/2007
    nom_de_famille: Rosso-Debord
    nom: Valérie Rosso-Debord
    type: depute
  depute_333421:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 333421
    extras:
      - conseil supérieur de la forêt, des produits forestiers et de la transformation du bois / membre titulaire
      - comité local d'information et de suivi du laboratoire souterrain de bure / membre titulaire
    adresses:
      - Permanence parlementaire 12 Rue Jean Errard 55000 Bar-le-Duc Téléphone : 03 29 70 69 76 Télécopie : 03 29 75 09 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 17 10 Télécopie : 01 40 63 17 11 
    circonscription: Meuse (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Pancher
    place_hemicycle: 326
    mails:
      - bpancher.depute@orange.fr
      - bpancher@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333421.asp
    profession: Directeur du développement
    site_web: http://www.bertrandpancher.com
    debut_mandat: 20/06/2007
    nom: Bertrand Pancher
    type: depute
  depute_333457:
    place_hemicycle: 143
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Premier vice-président de la Communauté de communes de la Côte des Mégalithes
      - Maire de Carnac, Morbihan (4444 habitants)
    sexe: H
    id_an: 333457
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333457.asp
    mails:
      - mgrall@assemblee-nationale.fr
      - michelgrall.depute@orange.fr
    adresses:
      - Permanence parlementaire 30 Avenue du Maréchal Foch 56400 Auray Téléphone : 02 97 56 24 24 Télécopie : 02 97 50 70 39 
      - Hôtel de ville BP 80 56341 Carnac Cedex Téléphone : 02 97 52 79 83 Télécopie : 02 97 52 79 78 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Morbihan (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Ingénieur conseil
    debut_mandat: 20/06/2007
    nom_de_famille: Grall
    nom: Michel Grall
    type: depute
  depute_333494:
    place_hemicycle: 494
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission de la défense nationale et des forces armées / membre / 
    sexe: F
    id_an: 333494
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333494.asp
    mails:
      - folivier@assemblee-nationale.fr
    adresses:
      - 21 Rue du Capitaine Lefort 56100 Lorient Téléphone : 02 97 21 26 63 Télécopie : 02 97 35 28 09 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Morbihan (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Chargée de mission auprès d'une collectivité territoriale
    debut_mandat: 20/06/2007
    nom_de_famille: Olivier-Coupeau
    nom: Françoise Olivier-Coupeau
    type: depute
  depute_333590:
    place_hemicycle: 57
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Saint-Avold, Moselle (16946 habitants)
    sexe: H
    id_an: 333590
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333590.asp
    mails:
      - wojciechowski1@orange.fr
      - awojciechowski@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 2 Boulevard de Lorraine 57500 Saint Avold Téléphone : 03 87 91 22 22 Télécopie : 03 87 91 14 63 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 62 27 Télécopie : 01 40 63 53 37 
    circonscription: Moselle (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Employé (secteur privé)
    debut_mandat: 20/06/2007
    nom_de_famille: Wojciechowski
    nom: André Wojciechowski
    type: depute
  depute_333611:
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 333611
    extras:
      - conseil d'administration de l'agence nationale pour l'amélioration des conditions de travail / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 93 17 
      - 11 Boulevard du Pont BP 7 57310 Guénange Téléphone : 03 82 50 70 20 
    circonscription: Moselle (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Filippetti
    place_hemicycle: 546
    mails:
      - afilippetti@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333611.asp
    profession: Enseignante et écrivain
    site_web: http://www.aureliefilippetti.org
    debut_mandat: 20/06/2007
    nom: Aurélie Filippetti
    type: depute
  depute_333818:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 333818
    adresses:
      - Mairie 59430 Saint-Pol-sur-Mer Téléphone : 03 28 29 66 00 Télécopie : 03 28 60 73 34 
      - Cabinet parlementaire 13 Rue Georges Pompidou 59279 Loor-Plage Téléphone : 03 28 63 09 54 Télécopie : 03 28 63 12 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (12ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Hutin
    place_hemicycle: 606
    autresmandats:
      - Maire de Saint-Pol-sur-Mer, Nord (23337 habitants)
      - Vice-président de la Communauté urbaine de Dunkerque
    mails:
      - hutinchristian@orange.fr
      - chutin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333818.asp
    profession: Médecin généraliste
    site_web: http://www.christianhutin.fr
    debut_mandat: 20/06/2007
    nom: Christian Hutin
    type: depute
  depute_333972:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: F
    id_an: 333972
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Espace Rive gauche (1er étage) 1 Avenue Jean Mabuse 59600 Maubeuge Téléphone : 03 27 62 35 32 Télécopie : 03 27 62 40 32 
    circonscription: Nord (23ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Marin
    place_hemicycle: 151
    autresmandats:
      - Membre du Conseil municipal de Jeumont, Nord (10775 habitants)
    mails:
      - christinemarin@orange.fr
      - cmarin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333972.asp
    profession: Commerçante
    site_web: http://www.christinemarin.fr
    debut_mandat: 20/06/2007
    nom: Christine Marin
    type: depute
  depute_333975:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 333975
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (24ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Pérat
    place_hemicycle: 627
    autresmandats:
      - Membre du conseil général (Nord)
      - Membre du Conseil municipal d'Anor, Nord (3093 habitants)
      - Premier vice-président de la Communauté de communes Action Fourmies et Environs
    mails:
      - jean-luc@perat.fr
      - jlperat@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/333975.asp
    profession: Professeur de l'enseignement secondaire et technique
    site_web: http://www.perat.fr
    debut_mandat: 20/06/2007
    nom: Jean-Luc Pérat
    type: depute
  depute_334116:
    place_hemicycle: 624
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Membre du conseil régional (Nord-Pas-de-Calais)
    sexe: F
    id_an: 334116
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334116.asp
    mails:
      - jmaquet@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 16 04 Télécopie : 01 40 63 16 06 
      - Permanence 10 Place Courbet 62000 Arras Téléphone : 03 21 24 66 49 Télécopie : 03 21 73 92 20 
    circonscription: Pas-de-Calais (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Directrice de mission
    debut_mandat: 20/06/2007
    nom_de_famille: Maquet
    nom: Jacqueline Maquet
    type: depute
  depute_334149:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 334149
    extras:
      - conseil national du littoral / membre titulaire
      - conseil national du tourisme / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Fasquelle
    place_hemicycle: 62
    autresmandats:
      - Maire du Touquet-Paris-Plage, Pas-de-Calais (5293 habitants)
      - Président de la Communauté de communes Mer et Terres d'Opale
    mails:
      - dfasquelle@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334149.asp
    profession: Professeur de faculté
    site_web: http://danielfasquelle.blogspot.com
    debut_mandat: 20/06/2007
    nom: Daniel Fasquelle
    type: depute
  depute_334160:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 334160
    adresses:
      - Mairie Place Godeffroy de Bouillon 62200 Boulogne sur Mer 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Cuvillier
    place_hemicycle: 371
    autresmandats:
      - Maire de Boulogne-sur-Mer, Pas-de-Calais (44862 habitants)
      - Président de la communauté d'agglomération du Boulonnais
    mails:
      - fcuvillier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334160.asp
    profession: Professeur de faculté
    site_web: http://www.fredericcuvillier.com
    debut_mandat: 20/06/2007
    nom: Frédéric Cuvillier
    type: depute
  depute_334525:
    place_hemicycle: 158
    fonctions:
      - commission des affaires culturelles et de l'éducation / secrétaire / 
    autresmandats:
      - Maire de Villeneuve-de-la-Raho, Pyrénées-Orientales (3625 habitants)
    sexe: F
    id_an: 334525
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334525.asp
    mails:
      - jirles@assemblee-nationale.fr
      - jacquelineirles@wanadoo.fr
    adresses:
      - Cabinet parlementaire 66180 Villeneuve de la Raho Téléphone : 04 68 56 76 38 Télécopie :  Télécopie : 04 68 87 11 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Orientales (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cadre supérieur
    debut_mandat: 20/06/2007
    nom_de_famille: Irles
    nom: Jacqueline Irles
    type: depute
  depute_334654:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 334654
    adresses:
      - Mairie 13 Rue Principale 68125 Houssen 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haut-Rhin (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Straumann
    place_hemicycle: 308
    autresmandats:
      - Membre du conseil général (Haut-Rhin)
      - Maire de Houssen, Haut-Rhin (1577 habitants)
    mails:
      - estraumann@assemblee-nationale.fr
      - ericstraumann@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334654.asp
    profession: Professeur agrégé
    site_web: http://www.ericstraumann.info
    debut_mandat: 20/06/2007
    nom: Éric Straumann
    type: depute
  depute_334750:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 334750
    adresses:
      - Permanence parlementaire 59 Ter Avenue du Point du Jour 69005 Lyon 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Havard
    place_hemicycle: 154
    autresmandats:
      - Membre du Conseil municipal de Lyon 5ème Arrondissement, Rhône (445523 habitants)
    mails:
      - mhavard@assemblee-nationale.fr
      - michel.havard.depute@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334750.asp
    profession: Autre cadre (secteur privé)
    site_web: http://www.michelhavard.fr
    debut_mandat: 20/06/2007
    nom: Michel Havard
    type: depute
  depute_334755:
    fonctions:
      - mision d'information commune sur la mesure des grandes données économiques et sociales / président / 
      - commission des finances / membre / 
    sexe: H
    id_an: 334755
    adresses:
      - 2 Place Louis Pradel 69001 Lyon 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Muet
    place_hemicycle: 549
    autresmandats:
      - Membre du Conseil municipal de Lyon 4ème Arrondissement, Rhône (445523 habitants)
    mails:
      - pamuet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334755.asp
    profession: Inspecteur général des finances
    site_web: http://pa-muet.com
    debut_mandat: 20/06/2007
    nom: Pierre-Alain Muet
    type: depute
  depute_334768:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 334768
    extras:
      - commision nationale d'agrément des associations représentant les usagers dans les instances hospitalières ou de santé publique / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 31 53 Téléphone : 01 40 63 31 03 Télécopie : 01 40 63 31 83 
      - Permanence parlementaire 117 Avenue de Saxe 69003 Lyon Téléphone : 04 37 45 49 49 Télécopie : 04 78 95 08 44 
    circonscription: Rhône (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Touraine
    place_hemicycle: 560
    autresmandats:
      - Membre de la communauté urbaine du Grand-Lyon
      - Adjoint au Maire de Lyon, Rhône (445523 habitants)
    mails:
      - jltouraine@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334768.asp
    profession: Professeur de médecine
    debut_mandat: 20/06/2007
    nom: Jean-Louis Touraine
    type: depute
  depute_334811:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / secrétaire / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 334811
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Télécopie : 01 40 63 31 97 
      - Permanence parlementaire 25 Rue Paul Verlaine 69100 Villeurbanne Téléphone : 04 78 84 09 12 Télécopie : 04 78 03 54 74 
    circonscription: Rhône (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Crozon
    place_hemicycle: 640
    autresmandats:
      - Membre du Conseil municipal de Villeurbanne, Rhône (124135 habitants)
    mails:
      - pcrozon@assemblee-nationale.fr
      - p.crozon@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334811.asp
    profession: Chargée de mission - Ancienne déléguée régionale chargée des droits des femmes
    site_web: http://blog.pascalecrozon.fr
    debut_mandat: 20/06/2007
    nom: Pascale Crozon
    type: depute
  depute_334843:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 334843
    adresses:
      - 1 Avenue Charles de Gaulle 69170 Tarare Téléphone : 04 74 05 29 59 Télécopie : 04 74 05 28 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Verchère
    place_hemicycle: 325
    autresmandats:
      - Maire de Cours-la-Ville, Rhône (4241 habitants)
    mails:
      - vercherepatrice@orange.fr
      - pverchere@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334843.asp
    profession: Assistant parlementaire
    site_web: http://www.patriceverchere.fr
    debut_mandat: 20/06/2007
    nom: Patrice Verchère
    type: depute
  depute_334906:
    place_hemicycle: 139
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Membre du Conseil municipal de Saint-Priest, Rhône (41023 habitants)
    sexe: H
    id_an: 334906
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334906.asp
    mails:
      - pmeunier@assemblee-nationale.fr
      - permanence.pmeunier@orange.fr
    adresses:
      - 18 Rue Louis Saunier 69330 Meyzieu Téléphone : 04 78 31 09 35 Télécopie : 04 78 31 72 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Rhône (13ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur de cabinet
    debut_mandat: 20/06/2007
    nom_de_famille: Meunier
    nom: Philippe Meunier
    type: depute
  depute_334951:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 334951
    adresses:
      - Permanence parlementaire 2 Rue Desault 70200 Lure Téléphone : 03 84 62 40 20 Télécopie : 03 84 62 40 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 15 78 Télécopie : 01 40 63 15 79 
    circonscription: Haute-Saône (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Jean-Michel Villaumé
    place_hemicycle: 567
    autresmandats:
      - Maire d'Héricourt, Haute-Saône (10129 habitants)
    mails:
      - permanence@depute-villaume.fr
      - jmvillaume@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334951.asp
    profession: Retraité de l'enseignement
    site_web: http://www.depute-villaume.fr
    debut_mandat: 20/06/2007
    nom: Jean-Michel Villaumé
    type: depute
  depute_334:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 334
    extras:
      - haut conseil de la coopération internationale / membre titulaire
    adresses:
      - Mairie 63114 Coudes Téléphone : 04 73 96 91 41 Télécopie : 04 73 96 69 63 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Puy-de-Dôme (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bacquet
    place_hemicycle: 411
    autresmandats:
      - Membre du conseil régional (Auvergne)
      - Maire de Coudes, Puy-de-Dôme (1109 habitants)
    mails:
      - jpbacquet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/334.asp
    profession: Médecin 
    debut_mandat: 20/06/2007
    nom: Jean-Paul Bacquet
    type: depute
  depute_335017:
    place_hemicycle: 405
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Président de la communauté d'agglomération de Chalon - Val de Bourgogne
      - Maire de Chalon-sur-Saône, Saône-et-Loire (50120 habitants)
    sexe: H
    id_an: 335017
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335017.asp
    mails:
      - csirugue@assemblee-nationale.fr
    adresses:
      - Permanence 22 Rue de la Banque 71100 Chalon-sur-Saône Téléphone : 03 85 90 04 30 Télécopie : 03 85 93 18 49 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Saône-et-Loire (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre supérieur (secteur privé)
    debut_mandat: 20/06/2007
    nom_de_famille: Sirugue
    nom: Christophe Sirugue
    type: depute
  depute_335040:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / vice-présidente / 
    sexe: F
    id_an: 335040
    adresses:
      - 111 Avenue Rhin et Danube 72000 Le Mans Téléphone : 02 43 28 32 33 Télécopie : 02 43 87 58 28 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Sarthe (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Labrette-Ménager
    place_hemicycle: 321
    autresmandats:
      - Membre du conseil général (Sarthe)
    mails:
      - fabienne.labrette.menagerlm1@orange.fr
      - flabrette@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335040.asp
    profession: Administrateur de sociétés
    site_web: http://www.fabienne-labrette-menager.com
    debut_mandat: 20/06/2007
    nom: Fabienne Labrette-Ménager
    type: depute
  depute_335054:
    fonctions:
      - commission des affaires européennes / secrétaire / 
      - mission d'information commune sur l'indemnisation des victimes des maladies nosocomiales et accès au dossier médical / membre / 
      - commission des lois / membre / 
    sexe: F
    id_an: 335054
    adresses:
      - Téléphone mobile : 06 31 65 46 63  contact@mariettakaramanli.fr
      - Permanence en circonscription 39 Rue Evrard  72100 Le Mans Téléphone : 02 43 86 91 91 Télécopie : 02 43 86 91 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Sarthe (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Karamanli
    place_hemicycle: 559
    autresmandats:
      - Adjointe au Maire du Mans, Sarthe (146105 habitants)
      - Membre de la Communauté Urbaine du Mans
    mails:
      - mkaramanli@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335054.asp
    profession: Professeur du secondaire et techn.
    site_web: http://www.mariettakaramanli.fr
    debut_mandat: 20/06/2007
    nom: Marietta Karamanli
    type: depute
  depute_335159:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 335159
    extras:
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre suppléant
    adresses:
      - 15, Avenue de Thônes 74000 Annecy Téléphone : 04 50 77 13 38 Télécopie : 04 50 77 19 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Savoie (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Tardy
    place_hemicycle: 157
    mails:
      - ltardy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335159.asp
    profession: Gérant d'entreprise
    site_web: http://tardy.hautetfort.com
    debut_mandat: 20/06/2007
    nom: Lionel Tardy
    type: depute
  depute_335319:
    place_hemicycle: 429
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 335319
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335319.asp
    mails:
      - smazetier@assemblee-nationale.fr
    adresses:
      - 263 Avenue Daumesnil 75012 Paris 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.sandrinemazetier.fr
    profession: Cadre supérieur (secteur privé)
    debut_mandat: 20/06/2007
    nom_de_famille: Mazetier
    nom: Sandrine Mazetier
    type: depute
  depute_335532:
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 335532
    adresses:
      - Permanence 8 Rue de la Cour des Noues 75020 Paris Téléphone : 01 43 15 61 24 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 64 Téléphone : 01 40 63 69 52 
    circonscription: Paris (21ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Pau-Langevin
    place_hemicycle: 451
    autresmandats:
      - Membre du Conseil municipal de Paris 20ème Arrondissement, Paris (182857 habitants)
    mails:
      - gpau@assemblee-nationale.fr
      - georgepaulangevin@yahoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335532.asp
    profession: Avocate
    site_web: http://www.georgepau-langevin.com
    debut_mandat: 20/06/2007
    nom: George Pau-Langevin
    type: depute
  depute_335543:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 335543
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 31 59 Télécopie : 01 40 63 31 89 
      - Permanence 23 Rue de la République 76100 Rouen  Téléphone : 02 77 76 47 55 Télécopie : 02 76 51 61 19 
    circonscription: Seine-Maritime (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Fourneyron
    place_hemicycle: 636
    autresmandats:
      - Maire de Rouen, Seine-Maritime (106512 habitants)
    mails:
      - vfourneyron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335543.asp
    profession: Médecin du sport
    site_web: http://www.valerie-fourneyron.parti-socialiste.fr
    debut_mandat: 20/06/2007
    nom: Valérie Fourneyron
    type: depute
  depute_335567:
    place_hemicycle: 153
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du Conseil municipal de Mont-Saint-Aignan, Seine-Maritime (21285 habitants)
    sexe: F
    id_an: 335567
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335567.asp
    mails:
      - fguegot@assemblee-nationale.fr
    adresses:
      - Autre téléphone : 02 22 51 01 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Maître de conférence associée
    debut_mandat: 20/06/2007
    nom_de_famille: Guégot
    nom: Françoise Guégot
    type: depute
  depute_335612:
    place_hemicycle: 577
    fonctions:
      - commission des affaires étrangères / secrétaire / 
    autresmandats:
      - Vice-président de la communauté de l'Agglomération Havraise
      - Maire de Gonfreville-l'Orcher, Seine-Maritime (9922 habitants)
    sexe: H
    id_an: 335612
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335612.asp
    mails:
      - jplecoq@assemblee-nationale.fr
      - jplecoq-6vgo@wanadoo.fr
    adresses:
      - Permanence 38 Rue des Marthyrs 76210 Bolbec Téléphone : 06 78 89 28 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (6ème)
    groupe:
      - gauche démocrate et républicaine / membre
    profession: Fonctionnaire de catégorie B
    debut_mandat: 20/06/2007
    nom_de_famille: Lecoq
    nom: Jean-Paul Lecoq
    type: depute
  depute_335758:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 335758
    extras:
      - commission nationale pour l'autonomie des jeunes / membre titulaire
    adresses:
      - Hôtel de ville 77120 Coulommiers Téléphone : 01 64 75 80 02 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-et-Marne (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Riester
    place_hemicycle: 224
    autresmandats:
      - Maire de Coulommiers, Seine-et-Marne (13852 habitants)
    mails:
      - friester@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335758.asp
    profession: Chef d'entreprise
    debut_mandat: 20/06/2007
    nom: Franck Riester
    type: depute
  depute_335999:
    place_hemicycle: 373
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 335999
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/335999.asp
    mails:
      - dbatho@assemblee-nationale.fr
    adresses:
      - Permanence de la Députée Place de la Mairie 79500 Melle Téléphone : 05 49 29 18 19 Télécopie : 05 49 29 11 33 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 94 16 
    circonscription: Deux-Sèvres (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre territorial
    debut_mandat: 20/06/2007
    nom_de_famille: Batho
    nom: Delphine Batho
    type: depute
  depute_336015:
    place_hemicycle: 372
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 336015
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336015.asp
    mails:
      - jgrellier@assemblee-nationale.fr
      - j.grellier@orange.fr
    adresses:
      - Permanence parlementaire 44 Rue Jean Jaurès 37 Résidence Démeter 79300 BRESSUIRE Téléphone : 05 49 74 58 38 Télécopie : 05 49 74 30 52 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Deux-Sèvres (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://jean-grellier.fr
    profession: Retraité salarié privé, dirigeant d'entreprise (SCOP)
    debut_mandat: 20/06/2007
    nom_de_famille: Grellier
    nom: Jean Grellier
    type: depute
  depute_336067:
    place_hemicycle: 478
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Vice-président du conseil général (Somme)
    sexe: H
    id_an: 336067
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336067.asp
    mails:
      - gilbert.mathon80@orange.fr
      - gmathon@assemblee-nationale.fr
    adresses:
      - Permanence 5 Rue du pont d'amour 80100 Abbeville Téléphone : 03 22 19 33 20 Télécopie : 03 22 19 12 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Somme (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Retraité de l'enseignement
    debut_mandat: 20/06/2007
    nom_de_famille: Mathon
    nom: Gilbert Mathon
    type: depute
  depute_336112:
    place_hemicycle: 573
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Vice-président du conseil général (Tarn)
    sexe: H
    id_an: 336112
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336112.asp
    mails:
      - jvalax@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 9 Avenue Kellermann-Cantepau 81000 Albi Téléphone : 05 63 80 29 25 Télécopie : 05 63 80 54 20 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Téléphone mobile : 06 70 51 37 61 
    circonscription: Tarn (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Valax
    nom: Jacques Valax
    type: depute
  depute_336175:
    place_hemicycle: 628
    fonctions:
      - commission des lois / membre / 
    sexe: F
    id_an: 336175
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336175.asp
    mails:
      - spinel@assemblee-nationale.fr
    adresses:
      - Permanence Parlementaire 71 Rue de l'Egalité 82100 Castelsarrasin Téléphone : 05 63 32 58 81 Télécopie : 05 63 32 09 95 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Tarn-et-Garonne (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    site_web: http://www.sylviapinel.com
    profession: Collaborateur de cabinet
    debut_mandat: 20/06/2007
    nom_de_famille: Pinel
    nom: Sylvia Pinel
    type: depute
  depute_336316:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 336316
    adresses:
      - 33, Cours Sadi Carnot BP 70044 84302 Cavaillon cedex Téléphone : 04 90 05 85 02 Télécopie : 04 90 71 29 58 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vaucluse (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bouchet
    place_hemicycle: 24
    autresmandats:
      - Maire de Cavaillon, Vaucluse (24497 habitants)
    mails:
      - jcbouchet@assemblee-nationale.fr
      - bouchetjc@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336316.asp
    profession: Gérant de société
    site_web: http://www.jeanclaudebouchet.fr
    debut_mandat: 20/06/2007
    nom: Jean-Claude Bouchet
    type: depute
  depute_336421:
    place_hemicycle: 611
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: F
    id_an: 336421
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336421.asp
    mails:
      - ccoutelle@assemblee-nationale.fr
    adresses:
      - 11 Place de France 86000 Poitiers Téléphone : 05 49 47 47 87 Télécopie : 05 49 47 47 86 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vienne (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.catherinecoutelle.fr
    profession: Retraitée de l'enseignement
    debut_mandat: 20/06/2007
    nom_de_famille: Coutelle
    nom: Catherine Coutelle
    type: depute
  depute_336439:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 336439
    adresses:
      - Permanence 1 Cité de la Roche BP 25 86160 Gençay Téléphone : 05 49 03 16 38 Télécopie : 05 49 03 16 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vienne (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Clément
    place_hemicycle: 612
    autresmandats:
      - Maire de Mauprévoir, Vienne (650 habitants)
    mails:
      - jmclement@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336439.asp
    profession: Avocat
    site_web: http://www.jeanmichelclement.com/
    debut_mandat: 20/06/2007
    nom: Jean-Michel Clément
    type: depute
  depute_336454:
    place_hemicycle: 610
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires culturelles et de l'éducation / secrétaire / 
    autresmandats:
      - Première adjointe de Limoges, Haute-Vienne (133907 habitants)
    sexe: F
    id_an: 336454
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336454.asp
    mails:
      - monique_boulestin@ville-limoges.fr
      - mboulestin@assemblee-nationale.fr
    adresses:
      - 40 Rue Haute Vienne 87000 Limoges Téléphone : 05 55 34 57 63 Télécopie : 05 55 34 38 83 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Vienne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur de lettres en détachement
    debut_mandat: 20/06/2007
    nom_de_famille: Boulestin
    nom: Monique Boulestin
    type: depute
  depute_336576:
    place_hemicycle: 230
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: F
    id_an: 336576
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336576.asp
    mails:
      - mlfort@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 36 Bis Rue de l'Epée 89100 Sens Téléphone : 03 86 65 47 83 Télécopie : 03 86 83 39 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yonne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.marielouisefort.fr
    debut_mandat: 20/06/2007
    nom_de_famille: Fort
    nom: Marie-Louise Fort
    type: depute
  depute_336898:
    fonctions:
      - commission des affaires culturelles et de l'éducation / secrétaire / 
    sexe: F
    id_an: 336898
    adresses:
      - Hôtel de Ville 57 Avenue Henri-Ravera 92220 Bagneux Téléphone : 01 46 65 49 00 Télécopie : 01 42 31 61 80 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 87 Télécopie : 01 40 63 54 63 
    circonscription: Hauts-de-Seine (11ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Amiable
    place_hemicycle: 580
    autresmandats:
      - Présidente de la Communauté d'agglomération Sud de Seine
      - Maire de Bagneux, Hauts-de-Seine (37225 habitants)
    mails:
      - mhamiable@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336898.asp
    profession: Enseignante
    site_web: http://www.mhamiable.fr
    debut_mandat: 20/06/2007
    nom: Marie-Hélène Amiable
    type: depute
  depute_336971:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 336971
    adresses:
      - Hôtel de ville 2 Rue de la Commune de Paris 93308 Aubervilliers cedex Téléphone : 01 48 39 52 39 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 93 26 Télécopie : 01 40 63 93 81 
    circonscription: Seine-Saint-Denis (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Goldberg
    place_hemicycle: 407
    autresmandats:
      - Membre du Conseil municipal de La Courneuve, Seine-Saint-Denis (34968 habitants)
    mails:
      - dgoldberg@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/336971.asp
    profession: Maître de conférences
    site_web: http://www.danielgoldberg.fr
    debut_mandat: 20/06/2007
    nom: Daniel Goldberg
    type: depute
  depute_337084:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 337084
    extras:
      - conseil de surveillance de la caisse nationale des allocations familiales / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 17 12 Télécopie : 01 40 63 17 14 
    circonscription: Seine-Saint-Denis (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gaudron
    place_hemicycle: 240
    autresmandats:
      - Membre du Conseil municipal d'Aulnay-sous-Bois, Seine-Saint-Denis (80018 habitants)
    mails:
      - ggaudron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337084.asp
    profession: Géologue
    site_web: http://ggaudron.fr
    debut_mandat: 20/06/2007
    nom: Gérard Gaudron
    type: depute
  depute_337171:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 337171
    extras:
      - conseil d'administration de l'établissement d'hospitalisation public de fresnes spécifiquement destine à l'accueil des personnes incarcérées / membre titulaire
    adresses:
      - Mairie Place de la vieille église 94290 Villeneuve-le-Roi Téléphone : 01 49 61 46 13 Télécopie : 01 45 97 39 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 23 
    circonscription: Val-de-Marne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Gonzales
    place_hemicycle: 152
    autresmandats:
      - Maire de Villeneuve-le-Roi, Val-de-Marne (18291 habitants)
    mails:
      - dgonzales@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337171.asp
    profession: Fonctionnaire
    site_web: http://www.didier-gonzales.fr
    debut_mandat: 20/06/2007
    nom: Didier Gonzales
    type: depute
  depute_337248:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 337248
    adresses:
      - Hôtel de ville Esplanade Georges Marrane 94200 Ivry Téléphone : 01.49.60.24.27 Télécopie : 01.72.04.64.89 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01.40.63.60.89 Télécopie : 01 40 63 61 92 
    circonscription: Val-de-Marne (10ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Gosnat
    place_hemicycle: 578
    autresmandats:
      - Maire d'Ivry-sur-Seine, Val-de-Marne (50908 habitants)
    mails:
      - pierregosnat@ivry94.fr
      - pgosnat@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337248.asp
    profession: Fonctionnaire
    site_web: http://www.pierregosnat.fr
    debut_mandat: 20/06/2007
    nom: Pierre Gosnat
    type: depute
  depute_337332:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 337332
    adresses:
      - Permanence 17 Avenue de l'Europe 95600 Eaubonne Téléphone : 01 39 59 73 10 Télécopie : 01 39 59 55 74 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 05 13 Télécopie : 01 40 63 05 93 
    circonscription: Val-d'Oise (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bodin
    place_hemicycle: 318
    autresmandats:
      - Membre du conseil régional (Ile-de-France)
    mails:
      - cbodin@assemblee-nationale.fr
      - bodin9504@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337332.asp
    profession: Attaché d'administration hospitalière
    site_web: http://www.claudebodin.fr
    debut_mandat: 20/06/2007
    nom: Claude Bodin
    type: depute
  depute_337421:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 337421
    adresses:
      - Permanence parlementaire 8 Rue de l'Hôtel Dieu 95500 Gonesse 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Paternotte
    place_hemicycle: 305
    autresmandats:
      - Maire de Sannois, Val-d'Oise (25353 habitants)
    mails:
      - abenard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337421.asp
    profession: Docteur en pharmacie, gérant de société pharmaceutique
    site_web: http://www.paternotte.fr
    debut_mandat: 20/06/2007
    nom: Yanick Paternotte
    type: depute
  depute_337442:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: F
    id_an: 337442
    adresses:
      - Immeuble "Le Negresco I" Boulevard Destrellau 97122 Baie Mahault Téléphone : 05 90 99 84 89 Télécopie : 05 90 99 73 88 
      - Mairie Boulevard des poissonniers 97126 Deshaies Téléphone : 05 90 28 57 09 Télécopie : 05 90 28 48 96 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 15 35 Téléphone : 01 40 63 15 36 Télécopie : 01 40 63 15 37 
    circonscription: Guadeloupe (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Marc
    place_hemicycle: 619
    autresmandats:
      - Maire de Deshaies, Guadeloupe (4039 habitants)
      - Membre de la Communauté de communes du Nord Basse Terre
    mails:
      - permanencejmarc@orange.fr
      - jmarc@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337442.asp
    profession: Retraité de l'enseignement
    site_web: http://www.jmlaguadeloupe.canalblog.com
    debut_mandat: 20/06/2007
    nom: Jeanny Marc
    type: depute
  depute_337483:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 337483
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 74 22 Téléphone : 01 40 63 74 23 Télécopie : 01 40 63 79 44 
    circonscription: Martinique (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Letchimy
    place_hemicycle: 409
    autresmandats:
      - Maire de Fort-de-France, Martinique (93986 habitants)
    mails:
      - sletchimy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337483.asp
    profession: Urbaniste
    site_web: http://serge-letchimy.fr
    debut_mandat: 20/06/2007
    nom: Serge Letchimy
    type: depute
  depute_337504:
    place_hemicycle: 629
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    autresmandats:
      - Vice-présidente du conseil régional (Guyane)
    sexe: F
    id_an: 337504
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337504.asp
    mails:
      - cberthelot@guyane.fr
      - cberthelot@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire PK 7 5 Route de Montjoly 97354 Remire Montjoly Téléphone : 05 94 25 02 96 Télécopie : 05 94 28 89 60 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Guyane (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    profession: Agricultrice
    debut_mandat: 20/06/2007
    nom_de_famille: Berthelot
    nom: Chantal Berthelot
    type: depute
  depute_337544:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 337544
    adresses:
      - Hôtel de ville 97430 Le Tampon 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 58 92 Télécopie : 01 40 63 99 04 
    circonscription: Réunion (3ème)
    groupe:
      - union pour un mouvement populaire / apparenté
    nom_de_famille: Robert
    place_hemicycle: 242
    autresmandats:
      - Maire du Tampon, Réunion (69849 habitants)
      - Président de la communauté de communes du Sud
    mails:
      - drobert@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337544.asp
    profession: Cadre administratif (collaborateur de cabinet)
    site_web: http://www.didierrobert.fr
    debut_mandat: 20/06/2007
    nom: Didier Robert
    type: depute
  depute_337550:
    place_hemicycle: 574
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire de Saint-Joseph, Réunion (30494 habitants)
    sexe: H
    id_an: 337550
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337550.asp
    mails:
      - plebreton@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Réunion (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Fonctionnaire de catégorie B
    debut_mandat: 20/06/2007
    nom_de_famille: Lebreton
    nom: Patrick Lebreton
    type: depute
  depute_337568:
    fonctions:
      - commission des affaires européennes / membre / 
      - mission d'information commune sur les prix des carburants dans les dom / membre / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 337568
    extras:
      - conseil supérieur de l'aviation marchande / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Réunion (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Fruteau
    place_hemicycle: 561
    autresmandats:
      - Maire de Saint-Benoît, Réunion (31662 habitants)
    mails:
      - jcfruteau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337568.asp
    profession: Retraité de l'enseignement
    debut_mandat: 20/06/2007
    nom: Jean-Claude Fruteau
    type: depute
  depute_337586:
    place_hemicycle: 73
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 337586
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337586.asp
    mails:
      - abdoulatifou.aly@orange.fr
      - aaly@assemblee-nationale.fr
    adresses:
      - 28  espace Coralium Route nationale 1 Kawéni,  BP 424 97600 Mamoudzou Téléphone : 02 69 61 18 71 Télécopie : 02 69 61 18 72 
      - 1  carrefour de la Liberté 97600 Mamoudzou 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Mayotte (1ère)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    profession: Avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Aly
    nom: Abdoulatifou Aly
    type: depute
  depute_337621:
    place_hemicycle: 323
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléant / 
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Papara, Polynésie Française (9659 habitants)
    sexe: H
    id_an: 337621
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337621.asp
    mails:
      - bsandras@assemblee-nationale.fr
      - bruno.sandras@papara.pf
    adresses:
      - Mairie 98712 Papara Téléphone : 00 689 54 75 47 Télécopie : 00 689 57 37 78 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Polynésie Française (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Permanent politique
    debut_mandat: 20/06/2007
    nom_de_famille: Sandras
    nom: Bruno Sandras
    type: depute
  depute_337633:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des finances / membre / 
    sexe: F
    id_an: 337633
    adresses:
      - 7 Rue René Autin BP 4477 97500 Saint-Pierre-et-Miquelon Téléphone : 05 08 41 99 98 Télécopie : 05 08 41 99 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 15 39 Télécopie : 01 40 63 15 40 
    circonscription: Saint-Pierre-et-Miquelon (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Girardin
    place_hemicycle: 621
    autresmandats:
      - Membre Conseil territorial de Saint-Pierre et Miquelon
    mails:
      - agirardin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337633.asp
    profession: Fonctionnaire de catégorie A
    site_web: http://www.annickgirardin.fr
    debut_mandat: 20/06/2007
    nom: Annick Girardin
    type: depute
  depute_337635:
    place_hemicycle: 558
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 337635
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/337635.asp
    mails:
      - alikuvalu@assemblee-nationale.fr
    adresses:
      - BP 82 98600 Mata Utu Téléphone : 00 681 72 26 02 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 16 34 
    circonscription: Wallis-et-Futuna (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    profession: Retraité de l'enseignement
    debut_mandat: 20/06/2007
    nom_de_famille: Likuvalu
    nom: Apeleto Albert Likuvalu
    type: depute
  depute_339:
    place_hemicycle: 626
    fonctions:
      - commission des finances / secrétaire / 
    autresmandats:
      - Premier vice-président de la communauté urbaine de Lille Métropole
      - Maire de Wattrelos, Nord (42764 habitants)
    sexe: H
    id_an: 339
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/339.asp
    mails:
      - dbaert@assemblee-nationale.fr
      - d.baert@ville-wattrelos.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Télécopie : 01 40 63 68 16 
      - Hôtel de Ville Place J. Delvainquière 59150 Wattrelos Téléphone : 03 20 81 64 97 
    circonscription: Nord (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Directeur à la Banque de France
    debut_mandat: 20/06/2007
    nom_de_famille: Baert
    nom: Dominique Baert
    type: depute
  depute_341339:
    place_hemicycle: 639
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du Conseil municipal de Thiviers, Dordogne (3261 habitants)
      - Membre du conseil général (Dordogne)
    sexe: F
    id_an: 341339
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/341339.asp
    circonscription: Dordogne (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Professeur
    debut_mandat: 07/03/2008
    nom_de_famille: Langlade
    nom: Colette Langlade
    type: depute
  depute_341481:
    place_hemicycle: 209
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 341481
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/341481.asp
    circonscription: Eure (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Médecin
    debut_mandat: 13/01/2009
    nom_de_famille: Lefrand
    nom: Guy Lefrand
    type: depute
  depute_341:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 341
    extras:
      - commission du dividende numérique / membre titulaire
    adresses:
      - Hôtel de Ville 26 Avenue André Morizet 92104 Boulogne-Billancourt Cedex Téléphone : 01 55 18 53 00 Télécopie : 01 55 18 63 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 60 00 Télécopie : 01 40 63 91 84 
    circonscription: Hauts-de-Seine (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Baguet
    place_hemicycle: 291
    autresmandats:
      - Maire de Boulogne-Billancourt, Hauts-de-Seine (105754 habitants)
    mails:
      - pc.baguet@mairie-boulogne-billancourt.fr
      - pcbaguet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/341.asp
    profession: Conseiller en communication
    site_web: http:// www.pcbaguet.com 
    debut_mandat: 20/06/2007
    nom: Pierre-Christophe Baguet
    type: depute
  depute_343034:
    place_hemicycle: 320
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Membre du conseil général (Maine-et-Loire)
      - Maire de Champigné, Maine-et-Loire (1896 habitants)
    sexe: H
    id_an: 343034
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/343034.asp
    circonscription: Maine-et-Loire (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Pharmacien d'officine
    debut_mandat: 20/07/2007
    nom_de_famille: Jeanneteau
    nom: Paul Jeanneteau
    type: depute
  depute_343385:
    place_hemicycle: 156
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire de Velaine-en-Haye, Meurthe-et-Moselle (1495 habitants)
    sexe: H
    id_an: 343385
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/343385.asp
    circonscription: Meurthe-et-Moselle (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chef d'entreprise
    debut_mandat: 20/04/2008
    nom_de_famille: Morenvillier
    nom: Philippe Morenvillier
    type: depute
  depute_343623:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des affaires sociales / membre / 
    autresmandats:
      - Membre du Conseil municipal de Roussy-le-Village, Moselle (962 habitants)
    sexe: F
    id_an: 343623
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/343623.asp
    circonscription: Moselle (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directrice des ventes
    debut_mandat: 17/11/2008
    nom_de_famille: Grommerch
    nom: Anne Grommerch
    type: depute
  depute_344878:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 344878
    adresses:
      - Permanence parlementaire 9 Rue Victor Hugo 69700 Givors Téléphone : 04 78 07 01 98 Télécopie : 04 72 24 00 09 
      - Permanence parlementaire 94 Boulevard des Allées 69420 Ampuis Téléphone : 04 74 56 90 77 Télécopie : 04 74 56 90 76 
      - Assemblée nationale 126 Rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 10 Télécopie : 01 40 63 56 70 
    circonscription: Rhône (11ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Durand
    place_hemicycle: 391
    autresmandats:
      - Maire de Chaponnay, Rhône (3317 habitants)
      - Vice-président du conseil général (Rhône)
    mails:
      - rdurand@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/344878.asp
    profession: Retraité
    site_web: http://www.raymond-durand.com
    debut_mandat: 02/06/2008
    nom: Raymond Durand
    type: depute
  depute_345727:
    place_hemicycle: 351
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Vice-président de la communauté d'agglomération Melun-Val-de-Seine
      - Maire de Melun, Seine-et-Marne (35591 habitants)
    sexe: H
    id_an: 345727
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/345727.asp
    circonscription: Seine-et-Marne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Proviseur-adjoint en retraite
    debut_mandat: 20/04/2008
    nom_de_famille: Millet
    nom: Gérard Millet
    type: depute
  depute_345898:
    place_hemicycle: 226
    fonctions:
      - commission des finances / membre / 
    sexe: F
    id_an: 345898
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/345898.asp
    circonscription: Yvelines (8ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 17/04/2009
    nom_de_famille: Dumoulin
    nom: Cécile Dumoulin
    type: depute
  depute_345937:
    place_hemicycle: 47
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Membre du Conseil municipal de Rambouillet, Yvelines (24758 habitants)
    sexe: H
    id_an: 345937
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/345937.asp
    circonscription: Yvelines (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chef d'entreprise
    debut_mandat: 20/07/2007
    nom_de_famille: Poisson
    nom: Jean-Frédéric Poisson
    type: depute
  depute_346652:
    place_hemicycle: 23
    fonctions:
      - commission des affaires sociales / membre / 
    autresmandats:
      - Maire d'Épinay-sur-Orge, Essonne (9399 habitants)
    sexe: H
    id_an: 346652
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/346652.asp
    circonscription: Essonne (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Administrateur civil hors classe
    debut_mandat: 20/07/2007
    nom_de_famille: Malherbe
    nom: Guy Malherbe
    type: depute
  depute_346692:
    place_hemicycle: 403
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: F
    id_an: 346692
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/346692.asp
    circonscription: Essonne (7ème)
    groupe:
      - union pour un mouvement populaire / apparenté
    profession: Ingénieur de recherche
    debut_mandat: 19/09/2008
    nom_de_famille: Briand
    nom: Françoise Briand
    type: depute
  depute_346886:
    place_hemicycle: 358
    fonctions:
      - commission des finances / membre / 
    autresmandats:
      - Membre du conseil régional (Ile-de-France)
    sexe: H
    id_an: 346886
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/346886.asp
    circonscription: Hauts-de-Seine (10ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/07/2007
    nom_de_famille: Lefebvre
    nom: Frédéric Lefebvre
    type: depute
  depute_346:
    place_hemicycle: 359
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Maire de Levallois-Perret, Hauts-de-Seine (54633 habitants)
    sexe: H
    id_an: 346
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/346.asp
    mails:
      - pbalkany@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence  43 Rue de Trebois 92300 Levallois-Perret Téléphone : 01 47 31 51 60 Télécopie : 01 47 37 49 47 
    circonscription: Hauts-de-Seine (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Directeur de société
    debut_mandat: 20/06/2007
    nom_de_famille: Balkany
    nom: Patrick Balkany
    type: depute
  depute_350:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 350
    extras:
      - comité consultatif de la législation et de la réglementation financières / membre suppléant
      - commission de surveillance de la caisse des dépôts et consignations / membre titulaire
    adresses:
      - Mairie 02140 Vervins Téléphone : 03 23 98 00 30 
      - Permanence 23 Rue du Général Leclerc 02140 Vervins Téléphone : 03 23 98 19 95 Télécopie : 03 23 98 15 00 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aisne (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Balligand
    place_hemicycle: 438
    autresmandats:
      - Maire de Vervins, Aisne (2653 habitants)
      - Membre du conseil général (Aisne)
    mails:
      - jp.balligand@wanadoo.fr
      - jpballigand@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/350.asp
    profession: Assistant parlementaire
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Balligand
    type: depute
  depute_356:
    fonctions:
      - commission des finances / membre / 
      - mission d'information commune sur les exonérations sociales / président / 
    sexe: H
    id_an: 356
    extras:
      - conseil de surveillance de la caisse nationale de l'assurance maladie des travailleurs salariés / membre titulaire
      - comité d'enquête sur le coût et le rendement des services publics / membre suppléant
      - comité de surveillance de la caisse d'amortissement de la dette sociale / membre titulaire
      - commission des comptes de la sécurité sociale / membre titulaire
    adresses:
      - 5 Rue Pierrette Louin Résidence L'Aiglon 31500 Toulouse Téléphone : 05 34 25 02 90 Télécopie : 05 34 25 02 99 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Hôtel de Ville 31240 Saint-Jean Téléphone : 05 61 37 63 02 Télécopie : 05 61 35 07 25 
    circonscription: Haute-Garonne (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bapt
    place_hemicycle: 437
    autresmandats:
      - Maire de Saint-Jean, Haute-Garonne (8362 habitants)
    mails:
      - depute.bapt@wanadoo.fr
      - gbapt@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/356.asp
    profession: Médecin cardiologue
    site_web: http://www.gerardbapt.info
    debut_mandat: 20/06/2007
    nom: Gérard Bapt
    type: depute
  depute_362:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 362
    extras:
      - conseil d'orientation de l'agence de la biomédecine / membre titulaire
    adresses:
      - Permanence 12 Place de la Halle 95220 Herblay Téléphone : 01 34 50 96 26 Télécopie : 01 34 50 94 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-d'Oise (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bardet
    place_hemicycle: 256
    autresmandats:
      - Membre du conseil régional (Ile-de-France)
    mails:
      - jbardet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/362.asp
    profession: Professeur de médecine
    debut_mandat: 20/06/2007
    nom: Jean Bardet
    type: depute
  depute_369:
    place_hemicycle: 174
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Troyes, Aube (60943 habitants)
      - Président de la communauté d'agglomération Troyenne (CAT)
    sexe: H
    id_an: 369
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/369.asp
    mails:
      - baroin.francois@wanadoo.fr
      - fbaroin@assemblee-nationale.fr
    adresses:
      - 33 Rue Urbain IV 10000 Troyes Téléphone : 03 25 73 09 70 Télécopie : 03 25 73 53 82 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Aube (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Avocat à la Cour
    debut_mandat: 20/06/2007
    nom_de_famille: Baroin
    nom: François Baroin
    type: depute
  depute_381:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 381
    adresses:
      - Hôtel du Département BP 193 93003 Bobigny Cedex 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (6ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bartolone
    place_hemicycle: 525
    autresmandats:
      - Président du conseil général (Seine-Saint-Denis)
    mails:
      - cbartolone@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/381.asp
    profession: Cadre de l'industrie pharmaceutique
    site_web: http://www.claudebartolone.net
    debut_mandat: 20/06/2007
    nom: Claude Bartolone
    type: depute
  depute_384:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 384
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Espace Soleil Route de Gruissan Bâtiment B, BP 134 11101 Narbonne cedex Téléphone : 04 68 90 28 28 Télécopie : 04 68 32 98 96 
    circonscription: Aude (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bascou
    place_hemicycle: 454
    autresmandats:
      - Président de la communauté d'agglomération de la Narbonnaise
      - Maire de Narbonne, Aude (51300 habitants)
    mails:
      - jbascou@assemblee-nationale.fr
      - permanence.bascou@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/384.asp
    profession: Cadre territorial
    site_web: http://www.jacques-bascou.fr
    debut_mandat: 20/06/2007
    nom: Jacques Bascou
    type: depute
  depute_390:
    place_hemicycle: 22
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du conseil régional (Basse Normandie)
    sexe: F
    id_an: 390
    extras:
      - conseil national de l'aménagement et du développement du territoire / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/390.asp
    mails:
      - sbassot@assemblee-nationale.fr
    adresses:
      - BP 20, Les Boëltières 61800 Le Ménil-Ciboult Téléphone : 02 33 66 60 20 Télécopie : 02 33 66 75 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Orne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Bassot
    nom: Sylvia Bassot
    type: depute
  depute_394:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 394
    adresses:
      - Secrétariat 26  Rue de Selle 59730 Solesmes Téléphone : 03 27 37 37 37 Télécopie : 03 27 37 38 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (22ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bataille
    place_hemicycle: 434
    autresmandats:
      - Membre du Conseil municipal de Solesmes, Nord (4767 habitants)
    mails:
      - cbataille@assemblee-nationale.fr
      - contact@christianbataille.org
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/394.asp
    profession: Professeur de lettres
    site_web: http://www.christianbataille.org
    debut_mandat: 20/06/2007
    nom: Christian Bataille
    type: depute
  depute_405480:
    place_hemicycle: 440
    fonctions:
      - commission des affaires économiques / membre / 
    autresmandats:
      - Maire de Sarcelles, Val-d'Oise (58002 habitants)
    sexe: H
    id_an: 405480
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/405480.asp
    mails:
      - fpupponi@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 Rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 57 Télécopie : 01 40 63 56 03 
      - Cabinet du Député-Maire 4 Place de Navarre 95200 Sarcelles Téléphone : 01 34 38 21 22 Télécopie : 01 39 90 27 10 
    circonscription: Val-d'Oise (8ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Directeur divisionnaire des Impôts
    debut_mandat: 16/12/2007
    nom_de_famille: Pupponi
    nom: François Pupponi
    type: depute
  depute_410:
    place_hemicycle: 70
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Membre du Conseil municipal de Pau, Pyrénées-Atlantiques (81000 habitants)
    sexe: H
    id_an: 410
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/410.asp
    mails:
      - f.bayrou@lesdemocrates.fr
      - fbayrou@assemblee-nationale.fr
    adresses:
      - MoDem 133 Bis Rue de l'Université 75007 Paris Téléphone : 01 53 59 20 00 
      - Permanence 34 Rue Henri Faisans 64000 Pau Téléphone : 05 59 30 61 91 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Atlantiques (2ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    profession: Professeur agrégé de lettres
    debut_mandat: 20/06/2007
    nom_de_famille: Bayrou
    nom: François Bayrou
    type: depute
  depute_412525:
    place_hemicycle: 72
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Vice-président du conseil général (Vendée)
    sexe: H
    id_an: 412525
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/412525.asp
    circonscription: Vendée (5ème)
    groupe:
      - députés n'appartenant à aucun groupe / membre
    profession: Conseiller des affaires étrangères hors classe (en détachement)
    debut_mandat: 13/04/2008
    nom_de_famille: Souchet
    nom: Dominique Souchet
    type: depute
  depute_414:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 414
    adresses:
      - Mairie 10 Place Charles Digeon 94160 Saint-Mandé Téléphone : 01 49 57 78 10 Télécopie : 01 49 57 78 09 
      - 271 Avenue de la République 94120 Fontenay-sous-Bois 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Beaudouin
    place_hemicycle: 233
    autresmandats:
      - Maire de Saint-Mandé, Val-de-Marne (19697 habitants)
    mails:
      - pbeaudouin@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/414.asp
    profession: Consultant en communication et relations publiques
    site_web: http://patrickbeaudouin.over-blog.com
    debut_mandat: 20/06/2007
    nom: Patrick Beaudouin
    type: depute
  depute_417099:
    place_hemicycle: 235
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 417099
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/417099.asp
    mails:
      - arobinet@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 Rue de l'Université 75355 Paris 07 SP 
      - Permanence 9 Place Royale 51100 Reims Téléphone : 03 26 97 00 37 Télécopie : 03 26 06 60 00 
    circonscription: Marne (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.arnaud-robinet.fr
    profession: Enseignant - Chercheur - Praticien hospitalier
    debut_mandat: 15/12/2008
    nom_de_famille: Robinet
    nom: Arnaud Robinet
    type: depute
  depute_418:
    place_hemicycle: 26
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Vice-président du conseil général (Charente-Maritime)
    sexe: H
    id_an: 418
    mails:
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/418.asp
    circonscription: Charente-Maritime (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chirurgien des hôpitaux
    debut_mandat: 20/07/2007
    nom_de_famille: Beaulieu
    nom: Jean-Claude Beaulieu
    type: depute
  depute_441:
    place_hemicycle: 597
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Maire de Saint-Paul, Réunion (88254 habitants)
    sexe: F
    id_an: 441
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/441.asp
    mails:
      - hbello@assemblee-nationale.fr
      - huguette.bello@wanadoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 19  Chaussée Royale BP 69 97862 Saint-Paul cedex Téléphone : 02 62 22 60 82 Télécopie : 02 62 45 57 07 
    circonscription: Réunion (2ème)
    groupe:
      - gauche démocrate et républicaine / membre
    profession: Directrice d'école maternelle
    debut_mandat: 20/06/2007
    nom_de_famille: Bello
    nom: Huguette Bello
    type: depute
  depute_475:
    place_hemicycle: 191
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Membre du conseil général (Loiret)
    sexe: H
    id_an: 475
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/475.asp
    mails:
      - jlbernard@assemblee-nationale.fr
      - jl.bernard.depute@wanadoo.fr
    adresses:
      - 38 Rue de la République 45000 Orléans Téléphone : 02 38 62 92 50 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loiret (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chirurgien retraité
    debut_mandat: 20/06/2007
    nom_de_famille: Bernard
    nom: Jean-Louis Bernard
    type: depute
  depute_479:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 479
    extras:
      - conseil supérieur des prestations sociales agricoles / membre titulaire
      - comité de surveillance de l'établissement de gestion du fonds de financement des prestations sociales des non-salariés agricoles / membre titulaire
      - commission du fonds national pour l'archéologie préventive / membre suppléant
    adresses:
      - Mairie 1 Route de la Bazouge de Cheméré 53480 Vaiges Téléphone : 02 43 66 57 64 
      - 58  Avenue Carnot 53200 Château-Gontier Téléphone : 02 43 07 25 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 12 Route de la Bazouge 53480 Vaiges Téléphone : 02 43 66 57 64 Télécopie : 02 43 66 57 72 
    circonscription: Mayenne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bernier
    place_hemicycle: 278
    autresmandats:
      - Membre de la communauté de communes d'Erve et Charnie
      - Maire de Vaiges, Mayenne (1071 habitants)
      - Membre du conseil général (Mayenne)
    mails:
      - mbernier@assemblee-nationale.fr
      - marc.bernier53@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/479.asp
    profession: Chirurgien-dentiste
    debut_mandat: 20/06/2007
    nom: Marc Bernier
    type: depute
  depute_493:
    place_hemicycle: 113
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 493
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/493.asp
    mails:
      - besselat.depute@wanadoo.fr
      - jybesselat@assemblee-nationale.fr
    adresses:
      - Permanence 32 Rue Jules Lecesne 76600 Le Havre Téléphone : 02 35 41 38 38 Télécopie : 02 35 42 05 49 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    site_web: http://www.jeanyvesbesselat.com
    debut_mandat: 20/06/2007
    nom_de_famille: Besselat
    nom: Jean-Yves Besselat
    type: depute
  depute_503:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 503
    extras:
      - commission de suivi du mémorandum d'accord signe le 26 novembre 1996 entre la france et la fédération de russie / membre suppléant
      - commission nationale pour l'éducation, la science et la culture ( unesco ) / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Conseil général 13 Rue Docteur Romieu 04000 Digne-les-Bains Téléphone : 04 92 30 04 04 Télécopie : 04 92 32 35 80 
    circonscription: Alpes-de-Haute-Provence (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bianco
    place_hemicycle: 415
    autresmandats:
      - Président du conseil général (Alpes-de-Haute-Provence)
    mails:
      - jlbianco@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/503.asp
    profession: Conseiller d'Etat
    site_web: http://www.jean-louis-bianco.com
    debut_mandat: 20/06/2007
    nom: Jean-Louis Bianco
    type: depute
  depute_508:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: F
    id_an: 508
    adresses:
      - Permanence 28 Avenue Grünberg 32100 Condom Téléphone : 05 62 68 09 55 Télécopie : 05 62 68 09 55 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gers (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Biémouret
    place_hemicycle: 637
    autresmandats:
      - Vice-présidente du conseil général (Gers)
    mails:
      - biemouret.gisele@orange.fr
      - gbiemouret@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/508.asp
    profession: Assistante parlementaire
    site_web: http://gisele-biemouret.over-blog.fr
    debut_mandat: 20/06/2007
    nom: Gisèle Biémouret
    type: depute
  depute_513:
    fonctions:
      - mission d'information commune sur les prix des carburants dans les dom / membre / 
      - commission du développement durable et de l'aménagement du territoire / vice-président / 
    sexe: H
    id_an: 513
    extras:
      - conseil d'administration de l'agence des aires marines protégées / membre titulaire
      - comité de l'initiative française pour les récifs coralliens / membre titulaire
      - conseil d'administration du conservatoire de l'espace littoral et des rivages lacustres / membre titulaire
    adresses:
      - 18 Rue de la Prévôté 80140 Oisemont Téléphone : 03 22 25 05 62 Télécopie : 03 22 25 89 30 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Somme (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bignon
    place_hemicycle: 106
    autresmandats:
      - Membre du conseil général (Somme)
    mails:
      - jbignon@assemblee-nationale.fr
      - jerome@bignon.info
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/513.asp
    profession: Avocat au Barreau de Paris
    site_web: http://www.bignon.info
    debut_mandat: 20/06/2007
    nom: Jérôme Bignon
    type: depute
  depute_522:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 522
    adresses:
      - Permanence 5 Rue du Parc 25300 Pontarlier Téléphone : 03 81 38 88 80 Télécopie : 03 81 38 86 27 
      - Hôtel de Ville BP 53095 25503 Morteau Téléphone : 03 81 68 56 56 Télécopie : 03 81 67 25 09 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Doubs (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Binetruy
    place_hemicycle: 1
    autresmandats:
      - Président de la communauté de communes du Val-de-Morteau
      - Adjoint au Maire de Morteau, Doubs (6372 habitants)
    mails:
      - jean-marie.binetruy@wanadoo.fr
      - jmbinetruy@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/522.asp
    profession: Enseignant
    site_web: http://jeanmariebinetruy.blogspirit.com/
    debut_mandat: 20/06/2007
    nom: Jean-Marie Binetruy
    type: depute
  depute_525:
    fonctions:
      - commission des affaires étrangères / membre / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    sexe: H
    id_an: 525
    extras:
      - institut de radioprotection et de sûreté nucléaire / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - BP 59 74103 Annemasse cedex Téléphone : 04 50 92 15 39 Télécopie : 04 50 92 60 40 
    circonscription: Haute-Savoie (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Birraux
    place_hemicycle: 270
    autresmandats:
      - Membre du conseil général (Haute-Savoie)
    mails:
      - deputebirraux@orange.fr
      - cbirraux@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/525.asp
    profession: Ingénieur
    site_web: http://www.claudebirraux.com
    debut_mandat: 20/06/2007
    nom: Claude Birraux
    type: depute
  depute_538:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 538
    extras:
      - conseil national de l'aménagement et du développement du territoire / membre titulaire
      - commission nationale de présélection des pôles d'excellence rurale / membre titulaire
      - observatoire des terrritoires / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence 9  Rue de la Gare 67700 Saverne Téléphone : 03 88 91 25 88 
    circonscription: Bas-Rhin (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Blessig
    place_hemicycle: 201
    autresmandats:
      - Maire de Saverne, Bas-Rhin (11201 habitants)
    mails:
      - eblessig@assemblee-nationale.fr
      - depute@blessig.org
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/538.asp
    profession: Avocat
    site_web: http://www.blessig.org
    debut_mandat: 20/06/2007
    nom: Émile Blessig
    type: depute
  depute_542:
    fonctions:
      - commission des lois / membre / 
    sexe: H
    id_an: 542
    extras:
      - commission nationale de l'admission exceptionnelle au séjour / membre suppléant
      - comité de suivi de l'agence française de l'adoption / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 41 Rue Bobillot 75013 Paris Téléphone : 01 45 89 88 63 Télécopie : 01 45 89 04 16 
    circonscription: Paris (10ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Blisko
    place_hemicycle: 547
    autresmandats:
      - Adjoint au Maire d'arrondissement de Paris (13ème Arrondissement), Paris (171523 habitants)
    mails:
      - sblisko@assemblee-nationale.fr
      - blisko@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/542.asp
    profession: Médecin
    site_web: http://www.blisko2007.typepad.fr
    debut_mandat: 20/06/2007
    nom: Serge Blisko
    type: depute
  depute_543:
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    sexe: H
    id_an: 543
    extras:
      - conseil d'administration du centre hospitalier national d'ophtalmologie des quinze-vingts / membre titulaire
      - haut conseil des musées de france / membre titulaire
    adresses:
      - 7 Rue François de Neufchâteau 75011 Paris 
      - Mairie 11 Place Léon Blum 75536 Paris cedex 11 Téléphone : 01 53 27 11 11 Télécopie : 01 53 27 10 54 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bloche
    place_hemicycle: 453
    autresmandats:
      - Conseiller de Paris, Paris (2121291 habitants)
      - Maire d'arrondissement de Paris (11ème Arrondissement), Paris (149074 habitants)
      - Conseiller de Paris
    mails:
      - p.bloche@wanadoo.fr
      - pbloche@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/543.asp
    profession: Directeur commercial
    site_web: http://www.patrickbloche.org
    debut_mandat: 20/06/2007
    nom: Patrick Bloche
    type: depute
  depute_546:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 546
    adresses:
      - Cabinet du 1er adjoint, Hôtel de ville Quai du port 13002 Marseille Téléphone : 04 91 55 35 90 Télécopie : 04 91 14 62 84 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bouches-du-Rhône (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Blum
    place_hemicycle: 112
    autresmandats:
      - Adjoint au Maire de Marseille, Bouches-du-Rhône (798021 habitants)
    mails:
      - rblum@mairie-marseille.fr
      - rblum@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/546.asp
    profession: Avocat
    site_web: http://www.roland-blum.com
    debut_mandat: 20/06/2007
    nom: Roland Blum
    type: depute
  depute_551:
    place_hemicycle: 592
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Président de la communauté d'agglomération de la Porte du Hainaut
      - Maire de Saint-Amand-les-Eaux, Nord (17170 habitants)
    sexe: H
    id_an: 551
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/551.asp
    mails:
      - abocquet@assemblee-nationale.fr
    adresses:
      - Mairie 65  Grand'Place 59230 Saint-Amand-les-Eaux Téléphone : 03 27 22 49 71 Téléphone : 03 27 22 48 47 Télécopie : 03 27 22 48 46 
      - BP 60026 59731 Saint-Amand-les-Eaux Téléphone : 03 27 27 86 40 Télécopie : 03 27 27 86 27 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (20ème)
    groupe:
      - gauche démocrate et républicaine / membre
    profession: Éducateur spécialisé
    debut_mandat: 20/06/2007
    nom_de_famille: Bocquet
    nom: Alain Bocquet
    type: depute
  depute_560:
    place_hemicycle: 360
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Maire de Saint-Yrieix-la-Perche, Haute-Vienne (7251 habitants)
      - Président de la communauté de communes du Pays de Saint-Yrieix
    sexe: H
    id_an: 560
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/560.asp
    mails:
      - dboisserie@assemblee-nationale.fr
    adresses:
      - Permanence 23 Place de la Nation BP 15 87500 Saint-Yrieix-la-Perche Téléphone : 05 55 75 07 07 Télécopie : 05 55 75 00 30 
      - Mairie 87500 Saint-Yrieix-la-Perche Téléphone : 05 55 08 88 57 Télécopie : 05 55 08 88 89 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Vienne (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Architecte
    debut_mandat: 20/06/2007
    nom_de_famille: Boisserie
    nom: Daniel Boisserie
    type: depute
  depute_580:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 580
    extras:
      - commission supérieure des sites, perspectives et paysages / membre titulaire
    adresses:
      - Mairie Place de l'Hôtel de Ville 17000 La Rochelle Téléphone : 05 46 28 18 06 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Charente-Maritime (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bono
    place_hemicycle: 456
    autresmandats:
      - Maire de La Rochelle, Charente-Maritime (76584 habitants)
    mails:
      - maxime.bono@ville-larochelle.fr
      - mbono@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/580.asp
    profession: Inspecteur des impôts
    site_web: http://maximebono.over-blog.com
    debut_mandat: 20/06/2007
    nom: Maxime Bono
    type: depute
  depute_599:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 599
    extras:
      - commission consultative du secret de la défense nationale / membre titulaire
    adresses:
      - 1 Rue de Toulouse 35000 Rennes Téléphone : 02 99 79 54 52 Télécopie : 02 99 78 10 92 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ille-et-Vilaine (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Boucheron
    place_hemicycle: 539
    autresmandats:
      - Membre du Conseil municipal de Rennes, Ille-et-Vilaine (205925 habitants)
    mails:
      - jmboucheron@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/599.asp
    profession: Assistant d'Université
    site_web: http://www.jmboucheron.fr
    debut_mandat: 20/06/2007
    nom: Jean-Michel Boucheron
    type: depute
  depute_621:
    fonctions:
      - commission des affaires européennes / membre / 
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 621
    extras:
      - haut conseil du secteur public / membre titulaire
      - conseil national de l'information statistique / membre suppléant
    adresses:
      - Hôtel de Ville BP19 76301 Sotteville-lès-Rouen cedex Téléphone : 02 35 72 08 19 Télécopie : 02 35 72 88 75 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Maritime (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Bourguignon
    place_hemicycle: 520
    autresmandats:
      - Maire de Sotteville-lès-Rouen, Seine-Maritime (29561 habitants)
    mails:
      - p.bourguignon@mairie-sotteville-les-rouen.fr
      - pbourguignon@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/621.asp
    profession: Sociologue urbaniste
    site_web: http://www.pierrebourguignon.net
    debut_mandat: 20/06/2007
    nom: Pierre Bourguignon
    type: depute
  depute_624:
    fonctions:
      - commission spéciale chargée de vérifier et d'apurer les comptes / vice-présidente / 
      - commission des affaires étrangères / membre / 
    sexe: F
    id_an: 624
    adresses:
      - 1 Rue Jacques Camille Paris BP 24 33030 Bordeaux cedex Téléphone : 05 56 29 07 29 Télécopie : 05 56 39 94 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Gironde (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bourragué
    place_hemicycle: 197
    autresmandats:
      - Membre du Conseil municipal de Bordeaux, Gironde (214633 habitants)
    mails:
      - chantal.bourrague@wanadoo.fr
      - cbourrague@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/624.asp
    profession: Cadre commercial
    site_web: http://www.chantal-bourrague.net
    debut_mandat: 20/06/2007
    nom: Chantal Bourragué
    type: depute
  depute_627:
    place_hemicycle: 441
    fonctions:
      - délégation chargée des activités internationales / membre / 
      - commission des affaires culturelles et de l'éducation / membre / 
      - délégation chargée de la communication et de la presse / membre / 
      - assemblée nationale / secrétaire / 01/10/2008
    sexe: F
    id_an: 627
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/627.asp
    mails:
      - dbousquet@assemblee-nationale.fr
      - bousquetsb@wanadoo.fr
    adresses:
      - Permanence 39 Avenue des Promenades BP 4633 22046 Saint-Brieuc cedex 2 Téléphone : 02 96 68 27 32 Télécopie : 02 96 68 25 93 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Côtes-d'Armor (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Chef d'établissement
    debut_mandat: 20/06/2007
    nom_de_famille: Bousquet
    nom: Danielle Bousquet
    type: depute
  depute_633:
    fonctions:
      - commission des finances / vice-président / 
    sexe: H
    id_an: 633
    extras:
      - conseil supérieur du service public ferroviaire / membre titulaire
      - conseil national pour le développement, l'aménagement et la protection de la montagne / membre titulaire
      - conseil d'orientation des finances publiques / membre titulaire
      - conseil d'administration du fonds pour le développement de l'intermodalité dans les transports / membre titulaire
      - commission de surveillance de la caisse des dépôts et consignations / membre titulaire
    adresses:
      - Secrétariat du Conseil général Château des Ducs de Savoie BP 1802 73018 Chambéry cedex Téléphone : 04 79 96 73 22 Télécopie : 04 79 62 29 31 
      - Permanence parlementaire 16  Place de la Sous-Préfecture BP 41 73302 Saint-Jean-de-Maurienne Téléphone : 04 79 59 93 96 Télécopie : 04 79 59 97 62 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Savoie (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bouvard
    place_hemicycle: 184
    autresmandats:
      - Vice-président du conseil général (Savoie)
    mails:
      - mbouvard@assemblee-nationale.fr
      - mbouvard@cg73.fr
      - mbouvard@icor.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/633.asp
    profession: Chargé de mission
    site_web: http://www.michelbouvard.com
    debut_mandat: 20/06/2007
    nom: Michel Bouvard
    type: depute
  depute_634:
    place_hemicycle: 250
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 634
    extras:
      - conseil d'orientation stratégique du fonds de solidarité prioritaire / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/634.asp
    mails:
      - loicbouvard-ploermel@wanadoo.fr
      - lbouvard@assemblee-nationale.fr
    adresses:
      - 8 Rue des Forges 56800 Ploërmel Téléphone : 02 97 74 05 47 Télécopie : 02 97 74 10 82 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 68 80 Télécopie : 01 40 63 98 11 
    circonscription: Morbihan (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Conseil en management
    debut_mandat: 20/06/2007
    nom_de_famille: Bouvard
    nom: Loïc Bouvard
    type: depute
  depute_653:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre titulaire / 
      - commission des lois / membre / 
    sexe: H
    id_an: 653
    extras:
      - conseil national de l'enseignement supérieur et de la recherche / membre suppléant
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 49 68 
      - 8 Passage de Jouy 93200 Saint-Denis Téléphone : 01 48 09 43 59 
      - CA Plaine Commune 21 Rue Jules Rimet 93200 Saint Denis Téléphone : 01 55 93 57 89 Téléphone : 01 48 22 08 63 
    circonscription: Seine-Saint-Denis (2ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Braouezec
    place_hemicycle: 585
    autresmandats:
      - Membre du Conseil municipal de Saint-Denis, Seine-Saint-Denis (85823 habitants)
      - Président de la communauté d'agglomération de Plaine Commune
    mails:
      - patrick.braouezec@plainecommune.com.fr
      - pbraouezec@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/653.asp
    profession: Instituteur
    debut_mandat: 20/06/2007
    nom: Patrick Braouezec
    type: depute
  depute_654:
    fonctions:
      - commission des finances / secrétaire / 
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
    sexe: H
    id_an: 654
    extras:
      - observatoire de la sécurité des cartes de paiement  / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (7ème)
    groupe:
      - gauche démocrate et républicaine / membre
    nom_de_famille: Brard
    place_hemicycle: 583
    autresmandats:
      - Membre du Conseil municipal de Montreuil, Seine-Saint-Denis (90588 habitants)
    mails:
      - jpbrard@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/654.asp
    profession: Instituteur
    site_web: http://www.depute-brard.org
    debut_mandat: 20/06/2007
    nom: Jean-Pierre Brard
    type: depute
  depute_667:
    place_hemicycle: 97
    fonctions:
      - délégation chargée des représentants d'intérêts / membre / 
      - délégation spéciale chargée de la question des groupes d'intérêt / membre / 
      - commission de la défense nationale et des forces armées / membre / 
      - assemblée nationale / questeur / 27/06/2007
      - délégation chargée de l'informatique et des nouvelles technologies / questeur, membre / 
      - délégation chargée des activités internationales / questeur, membre / 
    autresmandats:
      - Maire de Saint-Cyr-sur-Loire, Indre-et-Loire (16421 habitants)
    sexe: H
    id_an: 667
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/667.asp
    mails:
      - pbriand@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville BP 139 37541 Saint-Cyr cedex Téléphone : 02 47 42 80 02 Télécopie : 02 47 42 80 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Indre-et-Loire (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Chef d'entreprise et assureur
    debut_mandat: 20/06/2007
    nom_de_famille: Briand
    nom: Philippe Briand
    type: depute
  depute_680:
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 680
    extras:
      - commission du dividende numérique / membre titulaire
    adresses:
      - Les Portes de Crolles Rond-Point du Rafour 38927 Crolles Téléphone : 04 76 92 18 96 Télécopie : 04 76 92 18 98 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Brottes
    place_hemicycle: 519
    autresmandats:
      - Maire de Crolles, Isère (8260 habitants)
    mails:
      - francois.brottes@wanadoo.fr
      - fbrottes@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/680.asp
    profession: Directeur associé de société
    site_web: http://www.francois-brottes.com
    debut_mandat: 20/06/2007
    nom: François Brottes
    type: depute
  depute_689:
    place_hemicycle: 593
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
    autresmandats:
      - Membre du Conseil municipal du Blanc-Mesnil, Seine-Saint-Denis (46936 habitants)
    sexe: F
    id_an: 689
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/689.asp
    mails:
      - mgbuffet@assemblee-nationale.fr
    adresses:
      - 2  Rue Carnot 93240 Stains Téléphone : 01 42 35 71 97 Télécopie : 01 48 27 39 86 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Seine-Saint-Denis (4ème)
    groupe:
      - gauche démocrate et républicaine / membre
    profession: Employée
    debut_mandat: 20/06/2007
    nom_de_famille: Buffet
    nom: Marie-George Buffet
    type: depute
  depute_690:
    place_hemicycle: 110
    fonctions:
      - commission des lois / membre / 
    autresmandats:
      - Maire de Papeete, Polynésie Française (23535 habitants)
    sexe: H
    id_an: 690
    mails:
      - michel.buillard@mail.pf
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/690.asp
    circonscription: Polynésie Française (1ère)
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 75 73 Télécopie : 01 40 63 79 36 
      - Mairie BP 106 98713 Papeete Téléphone : 00 689 41 57 04 Télécopie : 00 689 45 46 36 
    groupe:
      - union pour un mouvement populaire / membre
    profession: Fonctionnaire
    debut_mandat: 20/06/2007
    nom_de_famille: Buillard
    nom: Michel Buillard
    type: depute
  depute_691:
    fonctions:
      - commission des affaires européennes / membre / 
      - mission d'information commune sur les exonérations sociales / rapporteur / 
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 691
    extras:
      - commission centrale de classement des débits de tabac / membre titulaire
      - conseil de surveillance du fonds de réserve pour les retraites / membre titulaire
      - conseil d'administration de l'office franco-allemand pour la jeunesse / membre titulaire
      - commission des comptes de la sécurité sociale / membre titulaire
      - haut conseil pour l'avenir de l'assurance maladie / membre titulaire
    adresses:
      - 7 Rue du Château 67380 Lingolsheim Téléphone : 03 88 10 31 40 Télécopie : 03 88 10 31 44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Bas-Rhin (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Bur
    place_hemicycle: 178
    autresmandats:
      - Maire de Lingolsheim, Bas-Rhin (16705 habitants)
    mails:
      - ybur@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/691.asp
    profession: Chirurgien-dentiste
    debut_mandat: 20/06/2007
    nom: Yves Bur
    type: depute
  depute_704:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / vice-président / 
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 704
    extras:
      - comité de gestion du fonds de soutien aux hydrocarbures ou assimiles d'origine nationale / membre titulaire
    adresses:
      - Communauté urbaine de Lille 1, Rue du Ballon BP 749 59000 Lille Téléphone : 03 20 21 22 23 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Nord (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Cacheux
    place_hemicycle: 625
    autresmandats:
      - Vice-président de la communauté urbaine de Lille Métropole
      - Membre du Conseil municipal de Lille, Nord (184231 habitants)
    mails:
      - acacheux@cudl-lille.fr
      - acacheux@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/704.asp
    profession: Ancien chargé d'études
    site_web: http://alain-cacheux.blogspirit.com/
    debut_mandat: 20/06/2007
    nom: Alain Cacheux
    type: depute
  depute_706:
    place_hemicycle: 536
    fonctions:
      - commission des finances / membre / 
      - mission d'information commune sur les prix des carburants dans les dom / rapporteur / 
    autresmandats:
      - Maire de Villeneuve-sur-Lot, Lot-et-Garonne (22772 habitants)
    sexe: H
    id_an: 706
    mails:
      - j.cahuzac@jcahuzac.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/706.asp
    circonscription: Lot-et-Garonne (3ème)
    adresses:
      - Mairie Boulevard de la République BP 317 47307 Villeneuve-sur-Lot Cedex Téléphone : 05 53 70 20 00 Télécopie : 05 53 70 34 57 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Chirurgien
    debut_mandat: 20/06/2007
    nom_de_famille: Cahuzac
    nom: Jérôme Cahuzac
    type: depute
  depute_707:
    place_hemicycle: 284
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 707
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/707.asp
    mails:
      - dcaillaud@assemblee-nationale.fr
      - permanence@dominique-caillaud.com
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 29 Rue La Bruyère BP 261 85007 La-Roche-sur-Yon cedex Téléphone : 02 51 37 82 15 Télécopie : 02 51 62 06 24 
    circonscription: Vendée (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Gérant de société
    debut_mandat: 20/06/2007
    nom_de_famille: Caillaud
    nom: Dominique Caillaud
    type: depute
  depute_716:
    fonctions:
      - commission des affaires européennes / membre / 
      - commission des lois / membre / 
    sexe: H
    id_an: 716
    extras:
      - conseil national des transports / membre suppléant
      - conseil national pour le développement, l'aménagement et la protection de la montagne / membre titulaire
    adresses:
      - 4 Quai Nobel 66000 Perpignan Téléphone : 04 68 35 61 49 Télécopie : 04 68 35 62 48 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pyrénées-Orientales (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Calvet
    place_hemicycle: 146
    autresmandats:
      - Maire du Soler, Pyrénées-Orientales (6862 habitants)
      - Vice-président de la Communauté d'agglomération Perpignan Méditerranée
    mails:
      - fcalvet@assemblee-nationale.fr
      - francois-calvet@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/716.asp
    profession: Avocat
    site_web: http://www.francois-calvet.com
    debut_mandat: 20/06/2007
    nom: François Calvet
    type: depute
  depute_719:
    place_hemicycle: 431
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 719
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/719.asp
    mails:
      - jccambadelis@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (20ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    site_web: http://www.cambadelis.net
    profession: Conseiller en communication
    debut_mandat: 20/06/2007
    nom_de_famille: Cambadélis
    nom: Jean-Christophe Cambadélis
    type: depute
  depute_732:
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / président / 
      - commission des finances / membre / 
    sexe: H
    id_an: 732
    adresses:
      - Hôtel de Ville 81500 Lavaur Téléphone : 05 63 83 12 20 Télécopie : 05 63 58 63 40 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Route de Castres Dominici 81500 Lavaur 
    circonscription: Tarn (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Carayon
    place_hemicycle: 348
    autresmandats:
      - Maire de Lavaur, Tarn (8537 habitants)
    mails:
      - boulzeb@yahoo.fr
      - bcarayon@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/732.asp
    profession: Avocat
    site_web: http://www.bcarayon-ie.com
    debut_mandat: 20/06/2007
    nom: Bernard Carayon
    type: depute
  depute_733:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 733
    extras:
      - commission supérieure du service public des postes et télécommunications / membre titulaire
    adresses:
      - Permanence parlementaire 34 Rue de l'Hôtel de Ville 81000 Albi Téléphone : 05 63 49 28 50 Télécopie : 05 63 49 28 54 
      - Conseil général Lices Georges Pompidou 81013 Albi cedex 9 Téléphone : 05 63 45 66 36 Télécopie : 05 63 45 64 43 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Tarn (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Carcenac
    place_hemicycle: 458
    autresmandats:
      - Président du conseil général (Tarn)
    mails:
      - tcarcenac@assemblee-nationale.fr
      - thierry.carcenac@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/733.asp
    profession: Inspecteur principal des impôts
    debut_mandat: 20/06/2007
    nom: Thierry Carcenac
    type: depute
  depute_734:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 734
    adresses:
      - 26 Rue de l'Abreuvoir 78570 Chanteloup-les-Vignes Téléphone : 01 39 70 88 99 Télécopie : 01 39 74 20 51 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Yvelines (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cardo
    place_hemicycle: 169
    autresmandats:
      - Président de la communauté de communes des Deux rives de la Seine
      - Membre du Conseil municipal de Chanteloup-les-Vignes, Yvelines (9544 habitants)
    mails:
      - caroline.raison@wanadoo.fr
      - pierre.cardo@wanadoo.fr
      - pcardo@assemblee-nationale.fr
      - claude.h.ney@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/734.asp
    profession: Cadre de gestion
    site_web: http://www.pierre-cardo.fr
    debut_mandat: 20/06/2007
    nom: Pierre Cardo
    type: depute
  depute_735:
    place_hemicycle: 448
    fonctions:
      - commission des affaires européennes / membre / 
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 735
    extras:
      - commission nationale de déontologie de la sécurité / membre titulaire
      - conseil d'orientation de l'observatoire national de la délinquance / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/735.asp
    mails:
      - caresche@club-internet.fr
      - ccaresche@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 76 Bis Rue Duhesme 75018 Paris Téléphone : 01 55 79 15 15 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Paris (18ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Chargé d'études
    debut_mandat: 20/06/2007
    nom_de_famille: Caresche
    nom: Christophe Caresche
    type: depute
  depute_746:
    place_hemicycle: 176
    fonctions:
      - commission des finances / rapporteur général / 
      - comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
      - commission des finances) de la mission d'évaluation et de contrôle (commission des finances) / (rapporteur général / 
    autresmandats:
      - Maire du Perreux-sur-Marne, Val-de-Marne (30057 habitants)
      - Membre de la Communauté d'agglomération de la Vallée de la Marne
    sexe: H
    id_an: 746
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/746.asp
    mails:
      - gcarrez@assemblee-nationale.fr
      - gillescarrez@leperreux.fr
    adresses:
      - Hôtel de Ville Place de la Libération 94170 Le Perreux-sur-Marne Téléphone : 01 48 71 53 53 Télécopie : 01 43 24 14 45 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Fonctionnaire de l'Etat en disponibilité
    debut_mandat: 20/06/2007
    nom_de_famille: Carrez
    nom: Gilles Carrez
    type: depute
  depute_765:
    place_hemicycle: 538
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    autresmandats:
      - Maire de Créteil, Val-de-Marne (82144 habitants)
    sexe: H
    id_an: 765
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/765.asp
    mails:
      - lcathala@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville 94000 Créteil Téléphone : 01 49 80 92 94 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Val-de-Marne (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Cadre hospitalier
    debut_mandat: 20/06/2007
    nom_de_famille: Cathala
    nom: Laurent Cathala
    type: depute
  depute_785:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - commission de la défense nationale et des forces armées / secrétaire / 
    sexe: H
    id_an: 785
    adresses:
      - Permanence parlementaire 9 Place de la République 50100 Cherbourg-Octeville 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Manche (5ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Cazeneuve
    place_hemicycle: 555
    autresmandats:
      - Maire de Cherbourg-Octeville, Manche (44108 habitants)
      - Président de la Communauté Urbaine de Cherbourg
    mails:
      - bcazeneuve@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/785.asp
    profession: Avocat au Barreau de Paris
    site_web: http://www.bernardcazeneuve.com
    debut_mandat: 20/06/2007
    nom: Bernard Cazeneuve
    type: depute
  depute_810:
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / membre / 
    sexe: H
    id_an: 810
    adresses:
      - Hôtel de Ville Place René Thimel 36300 Le Blanc Téléphone : 02 54 28 36 36 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - BP 107 36300 Le Blanc Téléphone : 02 54 37 18 30 Télécopie : 02 54 37 15 55 
    circonscription: Indre (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Chanteguet
    place_hemicycle: 461
    autresmandats:
      - Maire du Blanc, Indre (6997 habitants)
    mails:
      - jpchanteguet@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/810.asp
    profession: Conseiller économique
    site_web: http://chanteguet.com
    debut_mandat: 20/06/2007
    nom: Jean-Paul Chanteguet
    type: depute
  depute_815:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 815
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Permanence parlementaire 72 Rue de Paris 03200 Vichy Téléphone : 04 70 97 14 50 Télécopie : 04 70 97 00 26 
    circonscription: Allier (4ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / apparenté
    nom_de_famille: Charasse
    place_hemicycle: 614
    autresmandats:
      - Membre du conseil général (Allier)
    mails:
      - gcharasse@assemblee-nationale.fr
      - permanence.charasse@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/815.asp
    profession: Chargé de mission d'inspection de l'enseignement technique retraité
    site_web: http://www.charasse.net
    debut_mandat: 20/06/2007
    nom: Gérard Charasse
    type: depute
  depute_817:
    fonctions:
      - commission des affaires économiques / secrétaire / 
    sexe: H
    id_an: 817
    extras:
      - conseil de surveillance de l'agence de l'innovation industrielle / membre titulaire
      - conseil d'administration de l'établissement public de la cite des sciences et de l'industrie / membre titulaire
      - commission d'examen des pratiques commerciales / membre titulaire
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 69 23 Télécopie : 01 40 63 93 80 
      - 40  Mail ouest 45300 Pithiviers  Téléphone : 02 38 30 53 67 Télécopie : 02 38 30 15 74 
    circonscription: Loiret (5ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Jean-Paul Charié
    place_hemicycle: 248
    mails:
      - jpcharie@assemblee-nationale.fr
      - jean-paul.charie@orange.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/817.asp
    profession: Directeur multimédia de société de presse
    site_web: http://www.jeanpaulcharie.fr
    debut_mandat: 20/06/2007
    nom: Jean-Paul Charié
    type: depute
  depute_825:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 825
    adresses:
      - 250 Boulevard Saint-Germain 75007 Paris Téléphone : 01 42 22 69 51 Télécopie : 01 42 22 59 49 
      - Mairie 49410 Saint-Florent-le-Vieil Téléphone : 02 41 72 50 39 Télécopie : 02 41 72 55 85 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Maine-et-Loire (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Charette
    place_hemicycle: 193
    autresmandats:
      - Membre du conseil régional (Pays de la Loire)
      - Membre de la Communauté de communes du Canton de Saint-Florent-le-Vieil
      - Maire de Saint-Florent-le-Vieil, Maine-et-Loire (2623 habitants)
    mails:
      - hdecharette@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/825.asp
    profession: Avocat
    site_web: http://hervedecharette.typepad.fr
    debut_mandat: 20/06/2007
    nom: Hervé de Charette
    type: depute
  depute_856:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 856
    extras:
      - conseil national du bruit / membre suppléant
      - conseil d'orientation pour l'emploi / membre titulaire
    adresses:
      - Permanence 47 Rue de la Bolle 88100 Saint-Dié-des-Vosges Téléphone : 03 29 55 03 98 Télécopie : 03 29 55 07 61 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vosges (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cherpion
    place_hemicycle: 119
    autresmandats:
      - Membre du conseil régional (Lorraine)
    mails:
      - gcherpion@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/856.asp
    profession: Pharmacien
    debut_mandat: 20/06/2007
    nom: Gérard Cherpion
    type: depute
  depute_866:
    fonctions:
      - commission des affaires sociales / membre / 
    sexe: H
    id_an: 866
    extras:
      - conseil supérieur pour le reclassement professionnel et social des travailleurs handicapés / membre titulaire
      - conseil national consultatif des personnes handicapées / membre titulaire
      - conseil de la caisse nationale de solidarité pour l'autonomie / membre titulaire
    adresses:
      - 4 Rue Placette BP 141,  Moingt 42603 Montbrison cedex Téléphone : 04 77 58 37 36 Télécopie : 04 77 58 86 76 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Chossy
    place_hemicycle: 7
    autresmandats:
      - Membre du conseil régional (Rhône-Alpes)
    mails:
      - jfchossy@assemblee-nationale.fr
      - j-f.chossy@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/866.asp
    profession: Préparateur en pharmacie
    site_web: http://www.jeanfrancoischossy.fr
    debut_mandat: 20/06/2007
    nom: Jean-François Chossy
    type: depute
  depute_872:
    fonctions:
      - comité d'évaluation et de contrôle des politiques publiques / membre / 
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission des finances / membre / 
    sexe: H
    id_an: 872
    extras:
      - haut conseil des biotechnologies / membre suppléant
    adresses:
      - Hôtel de ville 86000 Poitiers Téléphone : 05 49 52 35 35 Télécopie : 05 49 41 91 97 
      - Permanence 16 Rue du Mouton 86000 Poitiers Téléphone : 05 49 50 97 79 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Vienne (1ère)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Claeys
    place_hemicycle: 426
    autresmandats:
      - Maire de Poitiers, Vienne (83448 habitants)
    mails:
      - aclaeys@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/872.asp
    profession: Enseignant
    debut_mandat: 20/06/2007
    nom: Alain Claeys
    type: depute
  depute_876:
    place_hemicycle: 249
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 876
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/876.asp
    mails:
      - pclement@assemblee-nationale.fr
    adresses:
      - Communauté de communes 42510 Balbigny 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire (6ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Avocat à la cour
    debut_mandat: 20/06/2007
    nom_de_famille: Clément
    nom: Pascal Clément
    type: depute
  depute_877:
    fonctions:
      - commission des affaires sociales / membre / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: F
    id_an: 877
    extras:
      - haut conseil de la famille / membre titulaire
      - conseil de surveillance de la caisse nationale des allocations familiales / membre titulaire
    adresses:
      - 11  Quai Turenne 44000 Nantes Téléphone : 02 40 35 74 74 Télécopie : 02 40 35 20 40 
      - Mairie Rue de l'Hôtel de ville 44000 Nantes Téléphone : 02 40 41 92 58 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Loire-Atlantique (2ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Clergeau
    place_hemicycle: 413
    autresmandats:
      - Adjointe au Maire de Nantes, Loire-Atlantique (269131 habitants)
      - Vice-présidente de la communauté urbaine de Nantes Métropole
    mails:
      - mfclergeau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/877.asp
    profession: Attachée commerciale
    site_web: http://www.clergeau.net
    debut_mandat: 20/06/2007
    nom: Marie-Françoise Clergeau
    type: depute
  depute_885:
    place_hemicycle: 600
    fonctions:
      - commission du développement durable et de l'aménagement du territoire / secrétaire / 
    sexe: H
    id_an: 885
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/885.asp
    mails:
      - ycochet@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 01 10 Télécopie : 01 40 63 01 90 
    circonscription: Paris (11ème)
    groupe:
      - gauche démocrate et républicaine / membre
    site_web: http://www.yvescochet.net
    profession: Informaticien
    debut_mandat: 20/06/2007
    nom_de_famille: Cochet
    nom: Yves Cochet
    type: depute
  depute_886:
    place_hemicycle: 632
    fonctions:
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Membre du Conseil municipal de Calais, Pas-de-Calais (77311 habitants)
    sexe: H
    id_an: 886
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/886.asp
    mails:
      - gcocquempot@assemblee-nationale.fr
    adresses:
      - Permanence parlementaire 64 Rue Berthois BP 473 62225 Calais cedex Téléphone : 03 21 19 11 20 Télécopie : 03 21 19 11 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Pas-de-Calais (7ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    profession: Chargé de mission
    debut_mandat: 20/06/2007
    nom_de_famille: Cocquempot
    nom: Gilles Cocquempot
    type: depute
  depute_891:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 891
    extras:
      - haut conseil du secteur public / membre titulaire
    adresses:
      - Permanence parlementaire 1  Rue Bonnat BP 14343 31028 Toulouse cedex 4 Téléphone : 05 61 14 00 31 Télécopie : 05 61 14 79 40 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Garonne (3ème)
    groupe:
      - socialiste, radical, citoyen et divers gauche / membre
    nom_de_famille: Cohen
    place_hemicycle: 542
    autresmandats:
      - Président de la communauté d'agglomération du Grand Toulouse
      - Maire de Toulouse, Haute-Garonne (390562 habitants)
    mails:
      - pcohen@assemblee-nationale.fr
      - contact@pierrecohen.net
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/891.asp
    profession: Ingénieur de recherche à l' INRIA
    site_web: http://www.pierrecohen.net
    debut_mandat: 20/06/2007
    nom: Pierre Cohen
    type: depute
  depute_909:
    fonctions:
      - commission des affaires sociales / secrétaire / 
      - mission d'évaluation et de contrôle des lois de financement de la sécurité sociale / membre / 
    sexe: H
    id_an: 909
    extras:
      - conseil d'administration de l'office national des anciens combattants et victimes de guerre / membre titulaire
    adresses:
      - Permanence parlementaire BP 21 38440 Saint-Jean-de-Bournay Téléphone : 04 74 59 76 76 Télécopie : 04 74 59 76 70 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Isère (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Colombier
    place_hemicycle: 347
    autresmandats:
      - Membre du conseil général (Isère)
    mails:
      - georges.colombier@orange.fr
      - gcolombier@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/909.asp
    profession: Salarié de l'industrie
    site_web: http://www.georges-colombier.fr
    debut_mandat: 20/06/2007
    nom: Georges Colombier
    type: depute
  depute_911:
    place_hemicycle: 210
    fonctions:
      - commission chargée de l'application de l'article 26 de la constitution / membre suppléante / 
      - commission des affaires étrangères / membre / 
    autresmandats:
      - Maire de Saint-Cyr-sous-Dourdan, Essonne (951 habitants)
    sexe: F
    id_an: 911
    extras:
      - conseil national de la sécurité routière / membre titulaire
      - observatoire national de la sécurité des établissements scolaires et d'enseignement supérieur / membre suppléante
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/911.asp
    mails:
      - gcolot@assemblee-nationale.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - Mairie 1 Route de Paris 91410 Saint-Cyr-sous-Dourdan Téléphone : 01 64 59 01 29 Télécopie : 01 64 59 12 31 
    circonscription: Essonne (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    debut_mandat: 20/06/2007
    nom_de_famille: Colot
    nom: Geneviève Colot
    type: depute
  depute_917:
    place_hemicycle: 99
    fonctions:
      - commission des affaires culturelles et de l'éducation / membre / 
      - bureau du comité d'évaluation et de contrôle des politiques publiques / membre de droit / 
    autresmandats:
      - Maire de Meaux, Seine-et-Marne (49421 habitants)
    sexe: H
    id_an: 917
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/917.asp
    mails:
      - jfcope@assemblee-nationale.fr
    adresses:
      - Hôtel de Ville 2 Place de l'Hôtel de Ville 77100 Meaux Téléphone : 01 60 09 97 00 Télécopie : 01 60 23 25 78 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP Téléphone : 01 40 63 63 77 Télécopie : 01 40 63 50 88 
    circonscription: Seine-et-Marne (6ème)
    groupe:
      - union pour un mouvement populaire / président
    profession: Administrateur civil et avocat
    debut_mandat: 20/06/2007
    nom_de_famille: Jean-François Copé
    nom: Jean-François Copé
    type: depute
  depute_923:
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 923
    extras:
      - conseil supérieur de la réserve militaire / membre titulaire
      - conseil supérieur de la participation / membre titulaire
    adresses:
      - 37 Bis Rue Maréchal de Lattre de Tassigny 52100 Saint-Dizier Téléphone : 03 25 05 61 09 Télécopie : 03 25 05 39 97 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Haute-Marne (2ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cornut-Gentille
    place_hemicycle: 94
    autresmandats:
      - Maire de Saint-Dizier, Haute-Marne (30896 habitants)
      - Président de la Communauté de communes de Saint-Dizier - Der et Perthois
    mails:
      - fcornut@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/923.asp
    profession: Cadre d'entreprise
    debut_mandat: 20/06/2007
    nom: François Cornut-Gentille
    type: depute
  depute_934:
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 934
    extras:
      - commission supérieure des sites, perspectives et paysages / membre titulaire
      - conseil supérieur de l' administration pénitentiaire / membre titulaire
    adresses:
      - Mairie Place Chateaubriand 35407 Saint-Malo Téléphone : 02 99 40 71 01 Télécopie : 02 99 40 71 21 
      - La Banneville Le Clos des Peupliers Saint-Ideuc 35400 Saint-Malo 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Ille-et-Vilaine (7ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Couanau
    place_hemicycle: 173
    autresmandats:
      - Maire de Saint-Malo, Ille-et-Vilaine (50654 habitants)
    mails:
      - rcouanau@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/934.asp
    profession: Inspecteur général de l'administration de l'Éducation nationale retraité
    debut_mandat: 20/06/2007
    nom: René Couanau
    type: depute
  depute_942:
    fonctions:
      - mission d'évaluation et de contrôle (commission des finances) / membre / 
      - commission spéciale chargée de vérifier et d'apurer les comptes / membre / 
      - commission des finances / vice-président / 
      - comité d'évaluation et de contrôle des politiques publiques / vice-président / 
    sexe: H
    id_an: 942
    extras:
      - conseil d'administration de l'établissement public de financement et de restructuration / membre titulaire
    adresses:
      - 38 Rue de la Petite-Sainte 51300 Vitry-le-François Téléphone : 03 26 73 29 70 Télécopie : 03 26 72 18 12 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Marne (5ème)
    groupe:
      - nouveau centre / membre
    nom_de_famille: Courson
    place_hemicycle: 375
    autresmandats:
      - Maire de Vanault-les-Dames, Marne (331 habitants)
      - Membre du conseil général (Marne)
      - Président de la communauté de communes des Côtes-de-Champagne
    mails:
      - charles.de-courson@wanadoo.fr
      - cdecourson@assemblee-nationale.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/942.asp
    profession: Magistrat à la Cour des comptes (conseiller référendaire)
    debut_mandat: 20/06/2007
    nom: Charles de Courson
    type: depute
  depute_946:
    fonctions:
      - commission des affaires étrangères / membre / 
    sexe: H
    id_an: 946
    extras:
      - conseil d'administration de l'agence française pour le développement international des entreprises (ubifrance) / membre titulaire
    adresses:
      - 8 Rue du Puits Notre-Dame 50200 Coutances Téléphone : 02 33 19 03 20 Télécopie : 02 33 19 03 21 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Manche (3ème)
    groupe:
      - union pour un mouvement populaire / membre
    nom_de_famille: Cousin
    place_hemicycle: 175
    mails:
      - acousin@assemblee-nationale.fr
      - cousin.alain@wanadoo.fr
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/946.asp
    profession: Agent général d'assurances
    site_web: http://www.alaincousin.fr
    debut_mandat: 20/06/2007
    nom: Alain Cousin
    type: depute
  depute_951:
    place_hemicycle: 171
    fonctions:
      - commission des affaires économiques / membre / 
    sexe: H
    id_an: 951
    extras:
      - commission supérieure des sites, perspectives et paysages / membre titulaire
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/951.asp
    mails:
      - couve.jean-michel@wanadoo.fr
      - jmcouve@assemblee-nationale.fr
    adresses:
      - 5  traverse des Lices 83990 Saint-Tropez Téléphone : 04 94 97 64 39 Télécopie : 04 94 43 99 44 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Var (4ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Cardiologue
    debut_mandat: 20/06/2007
    nom_de_famille: Couve
    nom: Jean-Michel Couve
    type: depute
  depute_966:
    place_hemicycle: 85
    fonctions:
      - commission de la défense nationale et des forces armées / membre / 
    sexe: H
    id_an: 966
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/966.asp
    mails:
      - hcuq@assemblee-nationale.fr
      - hcuq.perm@wanadoo.fr
    adresses:
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
      - 15 Avenue Charles de Gaulle BP 90067 78410 Aubergenville Cedex Téléphone : 01 30 91 19 50 Télécopie : 01 30 95 28 33 
    circonscription: Yvelines (9ème)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Ancien fonctionnaire du ministère de l'intérieur
    debut_mandat: 20/06/2007
    nom_de_famille: Cuq
    nom: Henri Cuq
    type: depute
  depute_998:
    place_hemicycle: 342
    fonctions:
      - commission des finances / membre / 
    sexe: H
    id_an: 998
    url_an: http://www.assembleenationale.fr/13/tribun/fiches_id/998.asp
    mails:
      - permanence.dassault@wanadoo.fr
      - odassault@assemblee-nationale.fr
    adresses:
      - Permanence 11 Bis Boulevard Amyot-d'Inville 60000 Beauvais Téléphone : 03 44 45 78 48 Télécopie : 03 44 48 54 49 
      - Assemblée nationale 126 rue de l'Université 75355 Paris 07 SP 
    circonscription: Oise (1ère)
    groupe:
      - union pour un mouvement populaire / membre
    profession: Président de sociétés
    debut_mandat: 20/06/2007
    nom_de_famille: Dassault
    nom: Olivier Dassault
    type: depute
